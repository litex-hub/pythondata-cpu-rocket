../Small24/TLBroadcastTracker_2.sv