../Small18/Queue_93.sv