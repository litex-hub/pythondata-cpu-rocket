../Medium82/TLXbar.sv