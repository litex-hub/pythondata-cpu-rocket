../Small18/Repeater_1.sv