../Small11/AXI4IdIndexer_1.sv