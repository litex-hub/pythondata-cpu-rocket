../Full84/TilePRCIDomain.sv