../Small11/Queue_15.sv