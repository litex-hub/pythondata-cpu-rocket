../Small88/TLBroadcastTracker_2.sv