../Small24/TilePRCIDomain.sv