../Medium22/TLXbar.sv