../Small42/TLBroadcastTracker_2.sv