../Small22/TLBuffer_2.sv