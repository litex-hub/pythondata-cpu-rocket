../Small11/AsyncResetRegVec_w8_i0.sv