../Small41/TLFIFOFixer_3.sv