../Full12/TLB_1.sv