../Small88/TLBroadcastTracker.sv