../Small21/TLMonitor_34.sv