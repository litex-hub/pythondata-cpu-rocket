../Small81/TLDebugModule.sv