../Small22/TLError_1.sv