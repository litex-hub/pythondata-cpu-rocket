../Small11/Repeater.sv