../Small84/ProbePicker.sv