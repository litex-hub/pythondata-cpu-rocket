../Small42/TLMonitor_45.sv