../Full11/HellaCacheArbiter.sv