../Medium11/RocketTile.sv