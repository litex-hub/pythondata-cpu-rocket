../Full11/BankedStore.sv