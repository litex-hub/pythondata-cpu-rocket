../Small14/TLMonitor_22.sv