../Small41/TLFIFOFixer_4.sv