../Small11/LevelGateway.sv