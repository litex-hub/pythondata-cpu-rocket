../Small24/TLBroadcastTracker_1.sv