../Small12/TLBuffer_4.sv