../Small24/TLBroadcast.sv