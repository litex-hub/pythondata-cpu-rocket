../Small81/AsyncQueueSink_2.sv