../Small11/TLBroadcastTracker.sv