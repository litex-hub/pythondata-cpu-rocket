../Small11/Queue_78.sv