../Small41/ProbePicker.sv