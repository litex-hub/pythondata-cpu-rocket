../Small42/TLFIFOFixer_3.sv