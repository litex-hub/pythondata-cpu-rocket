../Small11/ClockSinkDomain_1.sv