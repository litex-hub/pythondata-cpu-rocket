../Medium44/TLXbar.sv