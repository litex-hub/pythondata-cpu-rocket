../Small41/AXI4Buffer_1.sv