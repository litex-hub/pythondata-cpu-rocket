../Small41/TLBroadcastTracker.sv