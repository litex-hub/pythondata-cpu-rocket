../Small11/IntSyncAsyncCrossingSink_1.sv