../Small41/TLInterconnectCoupler_10.sv