../Small84/AXI4Buffer_1.sv