../Small11/Queue_73.sv