../Small22/TLBuffer_3.sv