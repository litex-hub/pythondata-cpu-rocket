../Linux11/DivSqrtRawFN_small_1.sv