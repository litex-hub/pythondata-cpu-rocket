../Medium12/SystemBus.sv