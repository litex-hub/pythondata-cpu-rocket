../Small11/ram_2x126.sv