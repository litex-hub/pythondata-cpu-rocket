../Medium41/Rocket.sv