../Linux11/FPToFP.sv