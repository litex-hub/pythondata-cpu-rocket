../Small41/Queue_48.sv