../Small81/TLInterconnectCoupler_17.sv