../Small11/TLBroadcastTracker_3.sv