../Small21/TLDebugModuleOuterAsync.sv