../Small44/BankBinder.sv