../Small81/TLMonitor_23.sv