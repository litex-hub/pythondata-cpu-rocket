../Medium41/TLPLIC.sv