../Small12/TLMonitor_23.sv