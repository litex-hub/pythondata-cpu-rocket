../Small22/TLMonitor_27.sv