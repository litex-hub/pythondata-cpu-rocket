../Small12/TLToAXI4_1.sv