../Small11/Queue_83.sv