../Medium81/TLPLIC.sv