../Linux11/RoundAnyRawFNToRecFN_2.sv