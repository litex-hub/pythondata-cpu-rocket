../Small11/PlusArgTimeout.sv