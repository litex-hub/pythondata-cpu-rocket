../Small81/TLMonitor_65.sv