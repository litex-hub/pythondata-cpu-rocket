../Small41/TLToAXI4_1.sv