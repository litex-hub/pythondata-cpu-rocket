../Medium12/TLMonitor_3.sv