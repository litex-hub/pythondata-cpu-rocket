../Small28/Queue_83.sv