../Full12/RocketTile.sv