../Small81/TLInterconnectCoupler_25.sv