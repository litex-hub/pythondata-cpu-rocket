../Small12/TLBuffer_2.sv