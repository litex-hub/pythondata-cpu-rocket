../Small11/DMIToTL.sv