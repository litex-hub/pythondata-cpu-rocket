../Small48/Queue_135.sv