../Small18/TLMonitor_21.sv