../Small21/Queue_45.sv