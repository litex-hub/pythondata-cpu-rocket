../Small11/mem_512x64.sv