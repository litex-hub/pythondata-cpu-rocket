../Small22/TLBuffer_4.sv