../Small11/OptimizationBarrier_22.sv