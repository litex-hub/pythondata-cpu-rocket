../Small42/TLMonitor_30.sv