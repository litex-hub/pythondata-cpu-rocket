../Small11/AsyncQueueSource.sv