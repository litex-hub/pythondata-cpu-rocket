../Small42/TLMonitor_32.sv