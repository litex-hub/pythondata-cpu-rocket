../Small42/TLXbar_16.sv