../Small41/AXI4UserYanker_1.sv