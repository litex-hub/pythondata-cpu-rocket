../Small21/TLBroadcastTracker.sv