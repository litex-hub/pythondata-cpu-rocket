../Small81/TLMonitor_35.sv