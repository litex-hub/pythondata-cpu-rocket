../Linux11/MulAddRecFNToRaw_preMul_1.sv