../Small41/TLMonitor_18.sv