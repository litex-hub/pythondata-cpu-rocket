../Full11/cc_banks_16384x64.sv