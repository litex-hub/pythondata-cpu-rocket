../Small21/BroadcastFilter.sv