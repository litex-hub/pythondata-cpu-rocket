../Small41/Queue_63.sv