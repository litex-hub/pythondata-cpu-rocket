../Small81/Queue_67.sv