../Small11/SimAXIMem_1.sv