../Small21/TLError_1.sv