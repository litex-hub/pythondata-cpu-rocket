../Small21/TLMonitor_33.sv