../Small42/TLBuffer_5.sv