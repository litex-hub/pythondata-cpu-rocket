../Small21/TLFIFOFixer_4.sv