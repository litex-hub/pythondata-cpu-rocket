../Small11/Arbiter.sv