../Full11/Repeater_4.sv