../Small11/TLInterconnectCoupler_11.sv