../Small11/NonSyncResetSynchronizerPrimitiveShiftReg_d3.sv