../Small42/TLMonitor_12.sv