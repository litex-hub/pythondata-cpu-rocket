../Small81/TLBuffer_5.sv