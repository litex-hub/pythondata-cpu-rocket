../Small42/TLMonitor_28.sv