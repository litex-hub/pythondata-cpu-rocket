../Small41/IntSyncCrossingSource_16.sv