../Small11/AsyncQueueSink_2.sv