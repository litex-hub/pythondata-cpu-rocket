../Small81/Repeater_3.sv