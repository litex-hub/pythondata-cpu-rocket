../Small11/TLDebugModuleInnerAsync.sv