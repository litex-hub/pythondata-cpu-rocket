../Small11/AsyncQueueSource_2.sv