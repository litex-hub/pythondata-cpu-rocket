../Small11/AsyncResetRegVec_w1_i0.sv