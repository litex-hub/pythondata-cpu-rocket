../Medium14/TLMonitor_1.sv