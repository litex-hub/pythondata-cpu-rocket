../Small12/TLXbar_10.sv