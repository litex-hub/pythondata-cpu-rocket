../Medium41/TLBuffer_10.sv