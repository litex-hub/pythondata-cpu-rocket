../Small24/BankBinder.sv