../Small82/TLFragmenter.sv