../Small22/TLMonitor_28.sv