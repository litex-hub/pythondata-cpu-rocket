../Small28/AXI4Fragmenter_1.sv