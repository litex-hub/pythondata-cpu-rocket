../Medium11/ShiftQueue.sv