../Small24/AXI4Xbar.sv