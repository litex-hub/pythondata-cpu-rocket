../Small81/TLMonitor_21.sv