../Linux11/IBuf.sv