../Small82/TLROM.sv