../Small21/MemoryBus.sv