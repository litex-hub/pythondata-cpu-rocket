../Medium44/TLMonitor_6.sv