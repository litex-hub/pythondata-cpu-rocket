../Small21/TLMonitor_16.sv