../Small82/TLBuffer_3.sv