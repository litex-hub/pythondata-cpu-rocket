../Small14/TLMonitor_23.sv