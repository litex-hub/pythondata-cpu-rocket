../Small11/ram_8x80.sv