../Small12/ProbePicker.sv