../Small11/TLFIFOFixer_2.sv