../Small22/TLBusBypassBar.sv