../Small12/TLROM.sv