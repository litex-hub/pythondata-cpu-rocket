../Small41/TLMonitor_25.sv