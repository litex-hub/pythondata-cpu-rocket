../Small14/TLMonitor_19.sv