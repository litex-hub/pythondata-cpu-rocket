../Small21/TLBuffer_4.sv