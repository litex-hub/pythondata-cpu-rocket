../Small14/Queue_72.sv