../Small81/IntXbar_9.sv