../Small22/TLError.sv