../Medium12/TLPLIC.sv