../Linux11/IntToFP.sv