../Small24/TLInterconnectCoupler_14.sv