../Medium44/TLBuffer_10.sv