../Small22/TLMonitor_22.sv