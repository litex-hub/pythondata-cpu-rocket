../Full11/ram_data_3x64.sv