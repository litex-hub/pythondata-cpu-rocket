../Small81/CSRFile.sv