../Small21/Queue_87.sv