../Medium11/TLXbar.sv