../Small81/Queue_15.sv