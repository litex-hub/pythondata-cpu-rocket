../Small22/TLAtomicAutomata_1.sv