../Small88/AXI4IdIndexer_2.sv