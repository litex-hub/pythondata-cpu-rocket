../Small82/TLFIFOFixer_2.sv