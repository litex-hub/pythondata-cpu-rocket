../Small11/Queue_40.sv