../Small82/TLMonitor_27.sv