../Small21/Queue_102.sv