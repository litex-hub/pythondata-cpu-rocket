../Small22/TLMonitor_35.sv