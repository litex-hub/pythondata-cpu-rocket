../Small44/AXI4Fragmenter_1.sv