../Small11/Queue_82.sv