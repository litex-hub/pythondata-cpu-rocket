../Small81/AXI4UserYanker.sv