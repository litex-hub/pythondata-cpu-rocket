../Small11/Queue_79.sv