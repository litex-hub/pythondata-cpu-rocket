../Medium14/SystemBus.sv