../Small21/TLMonitor_10.sv