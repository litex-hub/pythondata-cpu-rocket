../Small14/Repeater_1.sv