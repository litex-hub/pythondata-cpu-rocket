../Small88/Repeater_1.sv