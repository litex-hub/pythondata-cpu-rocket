../Medium22/TLMonitor_26.sv