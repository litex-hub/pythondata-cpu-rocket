../Small11/AXI4Fragmenter_2.sv