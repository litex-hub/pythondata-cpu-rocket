../Small82/ProbePicker.sv