../Small81/TLFragmenter_1.sv