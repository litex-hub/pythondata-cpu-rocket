../Small21/TLFIFOFixer_3.sv