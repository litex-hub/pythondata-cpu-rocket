../Small21/TLMonitor_17.sv