../Small12/TLWidthWidget_2.sv