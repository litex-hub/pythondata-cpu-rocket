../Small24/ProbePicker.sv