../Full11/Rocket.sv