../Small41/AsyncQueueSource_1.sv