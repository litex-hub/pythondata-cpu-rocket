../Small84/TLBroadcastTracker_2.sv