../Linux11/DivSqrtRawFN_small.sv