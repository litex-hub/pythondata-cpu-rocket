../Small11/TLMonitor.sv