../Medium84/TLMonitor_10.sv