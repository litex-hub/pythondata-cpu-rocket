../Small81/TLXbar_24.sv