../Small18/CoherenceManagerWrapper.sv