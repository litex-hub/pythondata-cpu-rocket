../Small11/AXI4ToTL.sv