../Medium84/TLFIFOFixer.sv