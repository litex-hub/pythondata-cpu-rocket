../Small21/TLMonitor_11.sv