../Small88/TLToAXI4_1.sv