../Small11/BankBinder.sv