../Small11/TLMonitor_26.sv