../Small11/TLBusBypass.sv