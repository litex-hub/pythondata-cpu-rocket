../Full11/RocketTile.sv