../Small11/TLMonitor_34.sv