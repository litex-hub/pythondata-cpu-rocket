../Linux11/CSRFile.sv