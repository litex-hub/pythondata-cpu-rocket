../Small81/Queue_159.sv