../Small82/Repeater_3.sv