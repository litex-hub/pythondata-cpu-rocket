../Small21/TLFragmenter_2.sv