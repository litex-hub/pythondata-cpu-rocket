../Linux11/Frontend.sv