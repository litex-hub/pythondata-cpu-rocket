../Small42/TLMonitor_27.sv