../Small88/AXI4Xbar.sv