../Small81/Queue_71.sv