../Small21/CLINT.sv