../Full11/head_21x6.sv