../Small81/TLFIFOFixer_4.sv