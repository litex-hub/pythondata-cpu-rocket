../Small24/TLMonitor_6.sv