../Small21/TLMonitor_21.sv