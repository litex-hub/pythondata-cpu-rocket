../Small28/TLInterconnectCoupler_2.sv