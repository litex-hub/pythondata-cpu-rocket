../Small84/Queue_105.sv