../Small21/AXI4Xbar.sv