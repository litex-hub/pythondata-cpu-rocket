../Small41/Queue_100.sv