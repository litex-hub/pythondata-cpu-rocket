../Medium11/IntSyncCrossingSource_8.sv