../Small21/IntSyncCrossingSource_8.sv