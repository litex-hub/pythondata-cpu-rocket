../Small22/CoherenceManagerWrapper.sv