../Small42/TLBuffer_2.sv