../Small48/MemoryBus.sv