../Small81/ram_9x11.sv