../Small84/TLInterconnectCoupler_2.sv