../Small42/TLMonitor_15.sv