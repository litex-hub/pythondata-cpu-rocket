../Small82/Queue_158.sv