../Small42/Queue_135.sv