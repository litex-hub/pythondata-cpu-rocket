../Small82/TLMonitor_29.sv