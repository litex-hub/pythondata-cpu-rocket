../Small88/Repeater.sv