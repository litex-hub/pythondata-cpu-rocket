../Small14/Queue_90.sv