../Small22/TLMonitor_7.sv