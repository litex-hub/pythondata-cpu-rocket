../Small11/TLMonitor_28.sv