../Small14/TLToAXI4_1.sv