../Small21/Queue_21.sv