../Small21/TLMonitor_15.sv