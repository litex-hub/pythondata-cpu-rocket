../Small88/TLInterconnectCoupler_26.sv