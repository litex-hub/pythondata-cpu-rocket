../Medium11/TLMonitor_1.sv