../Small28/TLBroadcastTracker_2.sv