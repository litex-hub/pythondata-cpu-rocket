../Small24/AXI4Buffer_1.sv