../Medium11/OptimizationBarrier.sv