../Medium42/ExampleRocketSystem.sv