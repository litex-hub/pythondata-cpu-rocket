../Small14/TLXbar.sv