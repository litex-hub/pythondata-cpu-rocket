../Small48/AXI4Xbar.sv