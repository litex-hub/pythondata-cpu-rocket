../Small21/TLMonitor_7.sv