../Small44/TLBroadcastTracker.sv