../Small81/Queue_37.sv