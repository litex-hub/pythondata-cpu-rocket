../Small48/TLInterconnectCoupler_18.sv