../Small22/TLMonitor_26.sv