../Small81/Queue_151.sv