../Linux11/DivSqrtRecFN_small_1.sv