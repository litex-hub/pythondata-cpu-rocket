../Small41/Queue_108.sv