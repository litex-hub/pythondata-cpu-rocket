../Small22/TLBroadcastTracker.sv