../Small11/TLBuffer_2.sv