../Small84/TLBroadcast.sv