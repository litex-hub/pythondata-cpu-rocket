../Small44/TLMonitor_25.sv