../Small12/TLMonitor_22.sv