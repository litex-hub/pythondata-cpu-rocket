../Small44/MemoryBus.sv