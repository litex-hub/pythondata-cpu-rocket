../Small11/Queue_34.sv