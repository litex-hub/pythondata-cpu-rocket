../Small41/TLMonitor_45.sv