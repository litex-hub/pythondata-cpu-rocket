../Medium42/SystemBus.sv