../Small81/AXI4Buffer_2.sv