../Small11/TLError_1.sv