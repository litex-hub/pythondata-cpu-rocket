../Small42/TLMonitor_19.sv