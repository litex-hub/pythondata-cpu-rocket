../Small22/TLMonitor_17.sv