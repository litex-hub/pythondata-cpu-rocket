../Small48/Queue_132.sv