../Medium82/TLBuffer_10.sv