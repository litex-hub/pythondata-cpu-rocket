../Small12/AXI4RAM.sv