../Medium81/TilePRCIDomain.sv