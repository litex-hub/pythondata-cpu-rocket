../Medium82/TLPLIC.sv