../Small82/TLMonitor_19.sv