../Small41/BroadcastFilter.sv