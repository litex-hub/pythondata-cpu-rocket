../Small21/TLMonitor_9.sv