../Small81/TLFragmenter_2.sv