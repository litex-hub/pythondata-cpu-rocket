../Small84/TLBroadcastTracker_3.sv