../Small21/TLMonitor_6.sv