../Small84/AXI4UserYanker_2.sv