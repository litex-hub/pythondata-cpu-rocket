../Full11/next_16x4.sv