../Small11/TLFragmenter_1.sv