../Small41/ClockCrossingReg_w21.sv