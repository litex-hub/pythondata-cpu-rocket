../Small84/TLBroadcastTracker.sv