../Small81/TLROM.sv