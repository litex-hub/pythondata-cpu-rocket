../Small81/TLToAXI4_1.sv