../Small11/ram_2x81.sv