../Small21/ClockSinkDomain.sv