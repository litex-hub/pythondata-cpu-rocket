../Small11/TLBusBypassBar.sv