../Small41/TLInterconnectCoupler_17.sv