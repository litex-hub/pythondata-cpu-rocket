../Small28/BankBinder.sv