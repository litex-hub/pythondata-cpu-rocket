../Small81/AXI4Fragmenter_1.sv