../Small12/TLBuffer_3.sv