../Medium81/CSRFile.sv