../Small81/PeripheryBus_1.sv