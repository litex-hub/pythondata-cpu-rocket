../Small21/TLInterconnectCoupler_13.sv