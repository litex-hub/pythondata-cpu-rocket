../Small22/BankBinder.sv