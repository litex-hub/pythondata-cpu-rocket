../Small21/TLToAXI4.sv