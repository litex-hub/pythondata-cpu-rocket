../Small82/TLMonitor_38.sv