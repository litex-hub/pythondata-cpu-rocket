../Small11/ram_2x6.sv