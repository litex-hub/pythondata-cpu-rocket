../Small41/Queue_109.sv