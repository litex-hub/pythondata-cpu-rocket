../Small41/TLMonitor_42.sv