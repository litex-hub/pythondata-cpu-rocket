../Small41/AXI4Xbar.sv