../Small41/TLMonitor_28.sv