../Small21/Queue_83.sv