../Small21/TLInterconnectCoupler_8.sv