../Small22/TLFragmenter.sv