../Small42/TLDebugModuleInner.sv