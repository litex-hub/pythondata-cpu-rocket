../Linux11/RoundAnyRawFNToRecFN_1.sv