../Small81/ProbePicker.sv