../Small28/TLBroadcastTracker.sv