../Small11/Queue_96.sv