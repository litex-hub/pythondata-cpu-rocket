../Small11/TLBuffer_3.sv