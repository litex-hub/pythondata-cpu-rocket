../Small81/TLBroadcastTracker.sv