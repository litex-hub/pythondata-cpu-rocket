../Small82/TLMonitor_70.sv