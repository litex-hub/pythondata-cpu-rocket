../Small21/CoherenceManagerWrapper.sv