../Small41/Queue_49.sv