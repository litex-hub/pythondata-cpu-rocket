../Small21/TLDebugModuleInnerAsync.sv