../Small12/TLFIFOFixer_3.sv