../Small21/TLMonitor_24.sv