../Small28/ProbePicker.sv