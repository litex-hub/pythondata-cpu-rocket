../Small48/Queue_129.sv