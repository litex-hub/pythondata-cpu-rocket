../Small81/TLMonitor_22.sv