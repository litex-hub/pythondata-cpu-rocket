../Small11/DCacheDataArray.sv