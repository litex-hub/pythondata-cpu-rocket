../Small81/TLXbar_5.sv