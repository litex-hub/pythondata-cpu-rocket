../Small41/PeripheryBus_1.sv