../Small12/TLMonitor_26.sv