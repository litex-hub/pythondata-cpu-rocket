../Small88/AXI4Fragmenter_1.sv