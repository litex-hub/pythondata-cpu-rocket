../Small48/TLMonitor_25.sv