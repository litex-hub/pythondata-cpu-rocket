../Small21/TLFragmenter.sv