../Small21/TLMonitor_14.sv