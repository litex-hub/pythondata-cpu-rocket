../Small24/Queue_83.sv