../Full11/TLB_1.sv