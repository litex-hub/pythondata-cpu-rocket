../Small41/TLInterconnectCoupler_13.sv