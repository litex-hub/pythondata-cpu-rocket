../Small24/TLMonitor_22.sv