../Small81/Queue_154.sv