../Small21/PeripheryBus_1.sv