../Small11/data_arrays_0_512x64.sv