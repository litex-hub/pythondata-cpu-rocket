../Small22/Queue_114.sv