../Small81/ram_2x82.sv