../Small21/BundleBridgeNexus_24.sv