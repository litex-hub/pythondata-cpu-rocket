../Small44/TLMonitor_10.sv