../Small81/TLMonitor_28.sv