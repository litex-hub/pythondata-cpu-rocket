../Small82/TLBroadcastTracker_2.sv