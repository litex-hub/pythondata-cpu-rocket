../Small22/TLROM.sv