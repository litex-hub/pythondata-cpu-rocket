../Linux11/RoundRawFNToRecFN.sv