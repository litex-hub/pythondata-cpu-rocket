../Small81/TLBroadcastTracker_2.sv