../Small12/TLInterconnectCoupler_12.sv