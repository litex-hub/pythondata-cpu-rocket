../Small11/AXI4Xbar_1.sv