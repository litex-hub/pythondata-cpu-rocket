../Small88/TLMonitor_37.sv