../Full11/next_40x6.sv