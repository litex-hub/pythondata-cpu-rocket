../Small11/OptimizationBarrier.sv