../Small44/TLFIFOFixer.sv