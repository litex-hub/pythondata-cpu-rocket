../Small11/AXI4Fragmenter.sv