../Small12/TLMonitor_12.sv