../Small41/TLROM.sv