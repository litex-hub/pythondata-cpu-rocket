../Small11/AXI4Xbar.sv