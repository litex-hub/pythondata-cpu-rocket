../Small81/TLMonitor_64.sv