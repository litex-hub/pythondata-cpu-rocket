../Linux11/RecFNToRecFN.sv