../Small18/TLMonitor_20.sv