../Small22/TLMonitor_40.sv