../Medium24/TLFIFOFixer.sv