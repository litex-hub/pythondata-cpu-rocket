../Medium11/Queue_78.sv