../Small24/TLToAXI4_1.sv