../Small24/TLFIFOFixer.sv