../Small81/Queue_70.sv