../Small44/ProbePicker.sv