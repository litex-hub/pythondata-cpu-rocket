../Medium22/TLFIFOFixer.sv