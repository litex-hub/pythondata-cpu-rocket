../Small22/TLMonitor_9.sv