../Medium42/TilePRCIDomain.sv