../Medium22/SystemBus.sv