../Small41/TLToAXI4.sv