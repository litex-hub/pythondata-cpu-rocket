../Small21/TLROM.sv