../Small24/TLMonitor_23.sv