../Small81/ClockCrossingReg_w29.sv