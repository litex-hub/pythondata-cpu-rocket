../Small42/TLBroadcastTracker_3.sv