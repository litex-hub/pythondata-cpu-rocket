../Small42/TLMonitor_26.sv