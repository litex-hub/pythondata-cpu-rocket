../Small21/TLBuffer_5.sv