../Small14/Queue_87.sv