../Small81/Queue_65.sv