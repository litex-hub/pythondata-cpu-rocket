../Small81/ram_2x11.sv