../Small21/Queue_98.sv