../Small14/TLBuffer_10.sv