../Small81/AXI4Fragmenter_2.sv