../Small12/TLMonitor_34.sv