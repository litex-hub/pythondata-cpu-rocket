../Linux11/regfile_32x65.sv