../Small22/TLAsyncCrossingSource.sv