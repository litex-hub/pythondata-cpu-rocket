../Small82/AXI4UserYanker_2.sv