../Small22/TLWidthWidget_2.sv