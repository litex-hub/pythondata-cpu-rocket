../Small42/TLFragmenter_3.sv