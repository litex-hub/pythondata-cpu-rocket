../Small48/TLMonitor_26.sv