../Full11/BreakpointUnit.sv