../Medium11/TLMonitor_24.sv