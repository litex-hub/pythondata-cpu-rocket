../Small81/Queue_60.sv