../Small11/TLBroadcastTracker_2.sv