../Small11/TLFragmenter_2.sv