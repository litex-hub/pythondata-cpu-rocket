../Small44/TLBroadcast.sv