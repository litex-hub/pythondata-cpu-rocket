../Small82/TLMonitor_34.sv