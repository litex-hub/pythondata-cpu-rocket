../Small21/Queue_89.sv