../Small11/Queue_5.sv