../Small28/AXI4Xbar.sv