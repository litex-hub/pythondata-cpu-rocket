../Small81/AXI4IdIndexer_2.sv