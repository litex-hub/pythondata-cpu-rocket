../Medium11/TLFIFOFixer.sv