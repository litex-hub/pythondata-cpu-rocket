../Small28/AXI4Buffer_1.sv