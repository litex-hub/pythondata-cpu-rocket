../Small42/AXI4Buffer_1.sv