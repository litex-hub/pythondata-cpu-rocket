../Small42/BankBinder.sv