../Medium11/TilePRCIDomain.sv