../Linux11/FPToInt.sv