../Small14/CoherenceManagerWrapper.sv