../Small11/TLMonitor_16.sv