../Small14/TLBroadcastTracker.sv