../Small81/TLMonitor_30.sv