../Linux11/INToRecFN.sv