../Small11/PeripheryBus_1.sv