../Small81/TLDebugModuleOuterAsync.sv