../Medium44/SystemBus.sv