../Medium14/TLBuffer_10.sv