../Small22/Queue_104.sv