../Small14/AXI4Buffer_1.sv