../Small41/TLBusBypassBar.sv