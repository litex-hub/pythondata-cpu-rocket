../Small81/TLBuffer_4.sv