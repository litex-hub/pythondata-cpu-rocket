../Small81/Queue_113.sv