../Small28/MemoryBus.sv