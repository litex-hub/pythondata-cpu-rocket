../Medium21/TLFIFOFixer.sv