../Small12/Repeater_4.sv