../Linux11/ShiftQueue.sv