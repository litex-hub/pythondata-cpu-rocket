../Small21/TLMonitor_35.sv