../Linux11/INToRecFN_1.sv