../Small41/Queue_128.sv