../Small82/Queue_168.sv