../Small28/TLWidthWidget_2.sv