../Small28/TLBroadcast.sv