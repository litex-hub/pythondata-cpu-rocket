../Small28/TLInterconnectCoupler_14.sv