../Small12/AXI4IdIndexer_2.sv