../Linux11/tag_array_64x84.sv