../Medium82/SystemBus.sv