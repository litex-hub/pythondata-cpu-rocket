../Small11/TLInterconnectCoupler_5.sv