../Small11/BundleBridgeNexus_15.sv