../Small11/TLFragmenter.sv