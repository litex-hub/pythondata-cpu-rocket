../Small12/Queue_100.sv