../Medium21/TLPLIC.sv