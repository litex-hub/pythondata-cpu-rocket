../Small82/TLMonitor_67.sv