../Small14/TLMonitor_4.sv