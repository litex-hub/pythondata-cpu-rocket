../Small82/TLXbar_24.sv