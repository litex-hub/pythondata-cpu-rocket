../Small12/TLAsyncCrossingSource.sv