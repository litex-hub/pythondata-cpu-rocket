../Small81/TLMonitor_68.sv