../Full82/RocketTile.sv