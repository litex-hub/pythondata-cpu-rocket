../Small11/tag_array_0_64x21.sv