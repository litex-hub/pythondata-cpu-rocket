../Small42/ProbePicker.sv