../Small41/AXI4IdIndexer.sv