../Small82/Queue_107.sv