../Full11/IDPool.sv