../Small82/TLMonitor_62.sv