../Medium44/TilePRCIDomain.sv