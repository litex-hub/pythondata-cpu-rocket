../Small41/TLMonitor_13.sv