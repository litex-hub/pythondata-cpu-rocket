../Small12/Repeater_3.sv