../Small82/TLMonitor_71.sv