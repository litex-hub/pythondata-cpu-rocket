../Small41/Queue_67.sv