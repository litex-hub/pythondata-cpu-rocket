../Small81/MemoryBus.sv