../Small28/TLBroadcastTracker_3.sv