../Small84/TLMonitor_36.sv