../Small81/TLMonitor_70.sv