../Small22/TLFragmenter_1.sv