../Small21/TLDebugModule.sv