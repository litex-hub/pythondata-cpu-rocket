../Small82/AXI4Xbar.sv