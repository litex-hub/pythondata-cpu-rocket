../Small14/BankBinder.sv