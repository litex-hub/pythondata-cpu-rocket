../Medium11/TLBuffer_10.sv