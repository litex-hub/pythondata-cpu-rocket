../Small41/TLInterconnectCoupler_11.sv