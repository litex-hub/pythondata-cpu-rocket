../Linux11/RecFNToIN.sv