../Full11/ram_2x111.sv