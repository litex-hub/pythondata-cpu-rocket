../Medium41/TLMonitor_6.sv