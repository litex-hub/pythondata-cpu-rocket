../Linux11/RecFNToIN_1.sv