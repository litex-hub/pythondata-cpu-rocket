../Small21/Queue_82.sv