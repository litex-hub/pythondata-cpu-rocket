../Full11/SinkA.sv