../Small11/CSRFile.sv