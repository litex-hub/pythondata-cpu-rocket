../Small21/AXI4Fragmenter_1.sv