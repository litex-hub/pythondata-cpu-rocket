../Small21/TLInterconnectCoupler_11.sv