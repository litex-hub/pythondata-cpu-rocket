../Small11/mem_268435456x64.sv