../Medium22/TLBuffer_10.sv