../Small11/TLMonitor_35.sv