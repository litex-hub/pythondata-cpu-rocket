../Small82/TLFragmenter_1.sv