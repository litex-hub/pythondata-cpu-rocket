../Small44/TilePRCIDomain.sv