../Full11/ListBuffer_2.sv