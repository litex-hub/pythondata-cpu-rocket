../Small12/TLInterconnectCoupler_2.sv