../Small12/TLMonitor_11.sv