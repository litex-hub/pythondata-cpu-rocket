../Small22/AXI4Xbar.sv