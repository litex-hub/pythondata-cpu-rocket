../Small11/TLMonitor_10.sv