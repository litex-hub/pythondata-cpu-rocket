../Small22/TLMonitor_20.sv