../Small81/TLMonitor_67.sv