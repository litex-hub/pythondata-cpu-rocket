../Small42/TLMonitor_46.sv