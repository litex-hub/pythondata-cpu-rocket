../Small12/AXI4Xbar.sv