../Small12/TLMonitor_4.sv