../Small18/AXI4Buffer_1.sv