../Small81/AXI4UserYanker_1.sv