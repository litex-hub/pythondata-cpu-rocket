../Small42/TLToAXI4.sv