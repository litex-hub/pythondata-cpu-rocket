../Small21/ClockCrossingReg_w17.sv