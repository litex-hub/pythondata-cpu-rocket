../Small41/Queue_106.sv