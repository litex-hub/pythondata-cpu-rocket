../Small14/Queue_93.sv