../Small81/TLToAXI4.sv