../Small84/TilePRCIDomain.sv