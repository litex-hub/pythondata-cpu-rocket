../Small82/TLAsyncCrossingSource.sv