../Linux11/DCacheDataArray.sv