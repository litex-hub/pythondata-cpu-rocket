../Linux11/CompareRecFN.sv