../Small11/TLMonitor_8.sv