../Small22/TLMonitor_14.sv