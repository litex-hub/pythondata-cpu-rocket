../Small41/TLMonitor_46.sv