../Small18/Repeater.sv