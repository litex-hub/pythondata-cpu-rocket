../Small41/CSRFile.sv