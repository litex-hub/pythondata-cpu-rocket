../Medium42/TLMonitor_31.sv