../Full44/TilePRCIDomain.sv