../Small88/MemoryBus.sv