../Small81/TLDebugModuleInnerAsync.sv