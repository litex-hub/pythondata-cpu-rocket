../Small82/TLMonitor_63.sv