../Small11/TLAsyncCrossingSource.sv