../Small12/TLMonitor_28.sv