../Small11/TLDebugModuleOuterAsync.sv