../Medium11/CSRFile.sv