../Small81/TLFragmenter_3.sv