../Small11/ram_4x8.sv