../Small88/Queue_107.sv