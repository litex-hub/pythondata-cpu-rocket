../Small81/TLInterconnectCoupler_26.sv