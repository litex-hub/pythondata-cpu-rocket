../Small81/IntSyncCrossingSource_32.sv