../Small12/TLBuffer_5.sv