../Small41/Rocket.sv