../Small81/TLMonitor_36.sv