../Small82/Repeater.sv