../Full11/ShiftQueue.sv