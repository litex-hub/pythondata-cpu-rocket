../Small41/Queue_130.sv