../Small14/Queue_74.sv