../Small42/AXI4Fragmenter_1.sv