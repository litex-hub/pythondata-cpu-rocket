../Small81/Queue_69.sv