../Small42/TLFragmenter_1.sv