../Small21/IntSyncCrossingSource_13.sv