../Small81/TLMonitor_31.sv