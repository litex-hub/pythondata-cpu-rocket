../Small41/TLBroadcastTracker_1.sv