../Small18/SimAXIMem.sv