../Small42/TLMonitor_42.sv