../Small21/FixedClockBroadcast.sv