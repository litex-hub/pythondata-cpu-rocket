../Small14/TilePRCIDomain.sv