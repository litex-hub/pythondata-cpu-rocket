../Small12/CLINT.sv