../Linux81/CSRFile.sv