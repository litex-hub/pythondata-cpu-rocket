../Medium24/TLBuffer_10.sv