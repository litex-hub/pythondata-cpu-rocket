../Small41/RocketTile.sv