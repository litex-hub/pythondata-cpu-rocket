../Small12/AXI4Buffer_2.sv