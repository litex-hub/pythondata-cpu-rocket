../Medium21/TLMonitor_27.sv