../Small21/TLMonitor_13.sv