../Small11/TLMonitor_33.sv