../Small12/TLMonitor_27.sv