../Small44/TLBroadcastTracker_3.sv