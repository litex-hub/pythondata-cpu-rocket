../Small21/AsyncQueueSink_2.sv