../Small81/TLMonitor_24.sv