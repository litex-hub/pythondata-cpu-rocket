../Linux11/RoundRawFNToRecFN_1.sv