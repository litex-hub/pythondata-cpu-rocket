../Small41/AXI4UserYanker_2.sv