../Medium24/TLMonitor_1.sv