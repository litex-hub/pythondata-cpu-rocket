../Linux11/DivSqrtRecFN_small.sv