../Small81/Queue_156.sv