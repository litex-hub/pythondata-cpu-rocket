../Small84/Queue_158.sv