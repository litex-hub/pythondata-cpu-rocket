../Medium81/TLMonitor_38.sv