../Small81/ram_2x117.sv