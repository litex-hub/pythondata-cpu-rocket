../Small14/Queue_80.sv