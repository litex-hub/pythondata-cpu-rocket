../Small11/FixedClockBroadcast.sv