../Small44/Queue_135.sv