../Linux11/DivSqrtRecFNToRaw_small_1.sv