../Small28/Queue_107.sv