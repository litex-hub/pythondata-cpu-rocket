../Small82/Queue_155.sv