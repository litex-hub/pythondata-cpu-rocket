../Medium21/TLXbar.sv