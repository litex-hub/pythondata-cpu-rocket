../Small11/TLMonitor_9.sv