../Linux11/MulAddRecFNPipe.sv