../Medium48/ExampleRocketSystem.sv