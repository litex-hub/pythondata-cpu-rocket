../Medium82/TLXbar_8.sv