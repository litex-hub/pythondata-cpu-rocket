../Small42/TLMonitor_16.sv