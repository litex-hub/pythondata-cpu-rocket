../Small12/TLBroadcast.sv