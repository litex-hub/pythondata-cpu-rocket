../Small12/TLMonitor_29.sv