../Small12/TLToAXI4.sv