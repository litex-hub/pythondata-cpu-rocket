../Full12/Frontend.sv