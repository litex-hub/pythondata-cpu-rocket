../Full11/Frontend.sv