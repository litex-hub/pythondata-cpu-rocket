../Medium14/TilePRCIDomain.sv