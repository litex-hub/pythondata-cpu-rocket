../Medium81/TLBuffer_10.sv