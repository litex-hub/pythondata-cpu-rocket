../Small81/ram_2x103.sv