../Small84/TLToAXI4_1.sv