../Small22/AXI4Buffer_1.sv