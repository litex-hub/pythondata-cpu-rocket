../Small11/TLInterconnectCoupler_7.sv