../Small11/TLFragmenter_3.sv