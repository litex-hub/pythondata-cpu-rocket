../Small11/RocketTile.sv