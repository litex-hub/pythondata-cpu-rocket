../Linux11/OptimizationBarrier_43.sv