../Small11/IntSyncSyncCrossingSink.sv