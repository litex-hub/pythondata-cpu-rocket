../Medium81/Queue_114.sv