../Small18/TLFIFOFixer_4.sv