../Small41/TLMonitor_11.sv