../Small41/TLFragmenter_2.sv