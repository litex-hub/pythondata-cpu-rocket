../Medium14/ExampleRocketSystem.sv