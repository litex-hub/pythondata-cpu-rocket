../Small41/AXI4Fragmenter_1.sv