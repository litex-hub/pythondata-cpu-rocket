../Small42/TLBuffer_3.sv