../Small22/Queue_83.sv