../Small82/TLXbar_8.sv