../Linux11/MulDiv.sv