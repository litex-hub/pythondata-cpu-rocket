../Small48/AXI4UserYanker_2.sv