../Small18/AXI4UserYanker_2.sv