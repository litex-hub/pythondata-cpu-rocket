../Small88/TLBroadcastTracker_3.sv