../Small41/Queue_62.sv