../Small82/TLMonitor_69.sv