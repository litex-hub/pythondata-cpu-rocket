../Medium12/TLMonitor_1.sv