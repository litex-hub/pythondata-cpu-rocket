../Small12/TLMonitor_18.sv