../Small81/TLMonitor_62.sv