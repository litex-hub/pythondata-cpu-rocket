../Medium82/TilePRCIDomain.sv