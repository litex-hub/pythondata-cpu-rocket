../Small11/TLMonitor_11.sv