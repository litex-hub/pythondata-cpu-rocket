../Small22/TLFragmenter_3.sv