../Medium24/TilePRCIDomain.sv