../Medium11/Queue_81.sv