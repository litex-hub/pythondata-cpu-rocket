../Small12/Queue_90.sv