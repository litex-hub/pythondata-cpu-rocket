../Small84/TLMonitor_35.sv