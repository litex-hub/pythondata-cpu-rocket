../Small42/Queue_101.sv