../Linux11/DCache.sv