../Small42/TLMonitor_13.sv