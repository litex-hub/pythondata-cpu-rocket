../Small12/TLMonitor_10.sv