../Small81/TLAtomicAutomata_1.sv