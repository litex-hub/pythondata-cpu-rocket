../Small42/TLMonitor_47.sv