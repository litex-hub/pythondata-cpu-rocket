../Small82/TLPLIC.sv