../Small81/ClockSinkDomain.sv