../Small84/TLMonitor_34.sv