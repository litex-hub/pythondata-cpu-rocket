../Small14/ram_2x264.sv