../Medium82/ExampleRocketSystem.sv