../Small11/PeripheryBus.sv