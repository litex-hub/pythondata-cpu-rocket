../Small82/TLMonitor_64.sv