../Linux11/RoundAnyRawFNToRecFN_3.sv