../Medium81/TLXbar_8.sv