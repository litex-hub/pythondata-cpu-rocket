../Small44/Queue_129.sv