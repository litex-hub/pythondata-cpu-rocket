../Small82/Repeater_4.sv