../Small81/Queue_13.sv