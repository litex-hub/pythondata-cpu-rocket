../Small11/ram_2x7.sv