../Small41/AXI4Buffer_2.sv