../Small18/TLBroadcastTracker_2.sv