../Small11/IntSyncCrossingSource_5.sv