../Small12/TLFIFOFixer_4.sv