../Medium11/HellaCacheArbiter.sv