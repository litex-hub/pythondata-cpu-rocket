../Small11/TLInterconnectCoupler_4.sv