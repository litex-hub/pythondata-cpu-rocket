../Small82/TLBuffer_4.sv