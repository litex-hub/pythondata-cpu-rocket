../Small12/TLMonitor_36.sv