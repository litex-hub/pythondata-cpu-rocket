../Small11/TLMonitor_32.sv