../Small84/AXI4Fragmenter_1.sv