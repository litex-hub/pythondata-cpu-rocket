../Small24/CoherenceManagerWrapper.sv