../Medium84/TLBuffer_10.sv