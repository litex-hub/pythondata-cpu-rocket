../Small81/AXI4Xbar.sv