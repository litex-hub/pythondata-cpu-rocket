../Small82/TLWidthWidget_2.sv