../Small88/TLMonitor_36.sv