../Small12/MemoryBus.sv