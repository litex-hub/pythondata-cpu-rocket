../Small11/PMPChecker.sv