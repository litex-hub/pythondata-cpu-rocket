../Small81/Queue_68.sv