../Small42/TLMonitor_48.sv