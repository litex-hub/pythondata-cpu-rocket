../Small11/SynchronizerShiftReg_w8_d3.sv