../Small81/TLFIFOFixer_3.sv