../Small41/TLMonitor_43.sv