../Small42/TLMonitor_44.sv