../Small22/TLMonitor_12.sv