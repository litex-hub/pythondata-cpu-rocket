../Small88/Queue_105.sv