../Small11/AsyncResetSynchronizerShiftReg_w1_d3_i0_1.sv