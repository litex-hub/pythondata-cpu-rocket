../Small42/TLMonitor_20.sv