../Small81/TLError_1.sv