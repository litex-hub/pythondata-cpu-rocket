../Small22/TLXbar_12.sv