../Small48/TLToAXI4_1.sv