../Small14/AXI4IdIndexer_2.sv