../Small81/AXI4IdIndexer.sv