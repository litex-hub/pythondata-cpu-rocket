../Medium11/Rocket.sv