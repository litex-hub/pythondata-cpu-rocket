../Full41/Rocket.sv