../Small11/ram_sink_2x2.sv