../Small24/TLInterconnectCoupler_2.sv