../Small82/AXI4Buffer_2.sv