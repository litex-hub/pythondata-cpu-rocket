../Small81/TLMonitor_33.sv