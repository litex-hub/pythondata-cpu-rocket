../Small42/CLINT.sv