../Small81/TLMonitor_9.sv