../Small11/TLFIFOFixer_3.sv