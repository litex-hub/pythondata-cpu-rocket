../Medium11/IBuf.sv