../Small14/AXI4RAM.sv