../Small82/TLAtomicAutomata_1.sv