../Small21/Queue_105.sv