../Small21/TLDebugModuleInner.sv