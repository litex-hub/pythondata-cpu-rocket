../Small28/TLBroadcastTracker_1.sv