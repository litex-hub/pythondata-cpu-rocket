../Small11/PLICFanIn.sv