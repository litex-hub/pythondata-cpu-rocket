../Small41/TLMonitor_27.sv