../Small41/Queue_9.sv