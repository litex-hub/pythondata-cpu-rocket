../Small88/TLBroadcast.sv