../Small21/TLMonitor_37.sv