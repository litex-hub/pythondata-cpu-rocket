../Small22/TLMonitor_39.sv