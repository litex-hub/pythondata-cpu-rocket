../Small81/Queue_158.sv