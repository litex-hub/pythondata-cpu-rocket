../Small88/TLBroadcastTracker_1.sv