../Small11/IntXbar_1.sv