../Medium14/TLXbar.sv