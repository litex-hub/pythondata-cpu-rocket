../Small18/AXI4RAM.sv