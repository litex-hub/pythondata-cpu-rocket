../Small82/Queue_161.sv