../Medium42/TLMonitor_32.sv