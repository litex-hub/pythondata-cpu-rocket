../Small42/AXI4UserYanker_2.sv