../Small11/IntXbar.sv