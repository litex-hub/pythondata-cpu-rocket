../Small11/TLXbar_10.sv