../Small21/AsyncQueueSource_1.sv