../Small81/Queue_106.sv