../Small22/TLMonitor_37.sv