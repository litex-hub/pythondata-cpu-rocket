../Small42/Queue_132.sv