../Small42/Queue_99.sv