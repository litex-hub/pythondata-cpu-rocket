../Medium22/TLMonitor_1.sv