../Small21/TLMonitor_40.sv