../Small81/TLInterconnectCoupler_11.sv