../Small24/Queue_89.sv