../Small12/TLXbar_8.sv