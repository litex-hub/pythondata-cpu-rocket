../Small21/AXI4UserYanker.sv