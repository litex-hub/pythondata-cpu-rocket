../Small12/AXI4UserYanker_2.sv