../Small12/TLError.sv