../Small11/TLMonitor_6.sv