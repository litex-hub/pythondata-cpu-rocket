../Small11/TLBroadcast.sv