../Small41/Queue_138.sv