../Small21/Queue_110.sv