../Small24/Queue_107.sv