../Small42/TLFIFOFixer_2.sv