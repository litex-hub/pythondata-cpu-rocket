../Medium11/Frontend.sv