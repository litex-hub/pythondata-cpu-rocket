../Small22/TLMonitor_16.sv