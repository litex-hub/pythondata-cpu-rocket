../Small41/TLBroadcastTracker_2.sv