../Linux41/Rocket.sv