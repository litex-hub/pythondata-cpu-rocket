../Small21/Queue_46.sv