../Small21/Queue_104.sv