../Small48/TLMonitor_29.sv