../Small22/TLMonitor_33.sv