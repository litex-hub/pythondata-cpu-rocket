../Small11/TLXbar_5.sv