../Small22/TLFIFOFixer_2.sv