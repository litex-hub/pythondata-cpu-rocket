../Small88/ProbePicker.sv