../Small14/TLInterconnectCoupler_2.sv