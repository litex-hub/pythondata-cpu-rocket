../Full11/data_16x65.sv