../Small88/TLWidthWidget_2.sv