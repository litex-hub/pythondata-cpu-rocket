../Small11/IntXbar_2.sv