../Small14/Repeater.sv