../Small81/Repeater_2.sv