../Medium11/PTW.sv