../Full11/Repeater.sv