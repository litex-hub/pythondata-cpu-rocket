../Small11/TLAtomicAutomata_1.sv