../Small11/AsyncResetRegVec_w2_i0.sv