../Medium12/TilePRCIDomain.sv