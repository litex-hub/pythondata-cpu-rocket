../Small84/TLFIFOFixer.sv