../Medium14/TLFIFOFixer.sv