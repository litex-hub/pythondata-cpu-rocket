../Small21/BankBinder.sv