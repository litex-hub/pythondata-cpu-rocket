../Small11/AXI4RAM.sv