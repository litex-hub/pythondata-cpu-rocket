../Small24/Queue_101.sv