../Small12/TLMonitor_32.sv