../Small28/TLToAXI4_1.sv