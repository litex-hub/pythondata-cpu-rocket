../Small11/ram_2x59.sv