../Small82/Repeater_1.sv