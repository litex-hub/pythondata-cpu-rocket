../Small11/TLMonitor_21.sv