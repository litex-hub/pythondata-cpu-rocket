../Small81/BankBinder.sv