../Small11/PMPChecker_2.sv