../Small82/TLMonitor_37.sv