../Small12/TLPLIC.sv