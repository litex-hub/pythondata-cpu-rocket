../Small24/TLBroadcastTracker_3.sv