../Small21/AXI4Fragmenter_2.sv