../Medium12/TLBuffer_10.sv