../Small14/TLFIFOFixer_4.sv