../Small42/TLToAXI4_1.sv