../Small88/TLMonitor_34.sv