../Small11/AsyncQueueSink_1.sv