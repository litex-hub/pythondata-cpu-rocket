../Small41/TLMonitor_16.sv