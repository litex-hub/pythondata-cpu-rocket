../Small18/TLBroadcastTracker.sv