../Small81/CLINT.sv