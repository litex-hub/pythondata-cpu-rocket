../Small21/Queue_31.sv