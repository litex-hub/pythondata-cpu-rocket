../Small21/TLFIFOFixer_2.sv