../Small21/Queue_49.sv