../Small42/TLPLIC.sv