../Small11/Queue_28.sv