../Small12/TLBroadcastTracker_2.sv