../Small42/TLInterconnectCoupler_18.sv