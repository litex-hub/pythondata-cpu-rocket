../Small12/TLMonitor_21.sv