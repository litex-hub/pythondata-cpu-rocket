../Small11/IBuf.sv