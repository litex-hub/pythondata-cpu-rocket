../Small41/TLMonitor_26.sv