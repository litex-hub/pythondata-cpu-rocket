../Small21/TLMonitor_18.sv