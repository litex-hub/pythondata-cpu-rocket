../Small21/AXI4Xbar_1.sv