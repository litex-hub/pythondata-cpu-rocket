../Full11/DCache.sv