../Small21/TLMonitor_8.sv