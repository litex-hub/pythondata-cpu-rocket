../Small42/TLAtomicAutomata_1.sv