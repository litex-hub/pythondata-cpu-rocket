../Small44/TLToAXI4_1.sv