../Small12/Queue_74.sv