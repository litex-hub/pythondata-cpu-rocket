../Small12/ram_4x144.sv