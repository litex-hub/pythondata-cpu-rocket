../Small12/TLBroadcastTracker_3.sv