../Small22/TLMonitor_10.sv