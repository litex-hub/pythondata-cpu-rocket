../Small22/ProbePicker.sv