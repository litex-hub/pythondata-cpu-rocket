../Linux11/OptimizationBarrier_42.sv