../Small11/Queue_27.sv