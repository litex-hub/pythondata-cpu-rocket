../Small11/OptimizationBarrier_21.sv