../Small84/TLInterconnectCoupler_26.sv