../Small81/CoherenceManagerWrapper.sv