../Full11/Arbiter.sv