../Small14/TLBroadcast.sv