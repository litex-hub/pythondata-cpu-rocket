../Small41/Queue_133.sv