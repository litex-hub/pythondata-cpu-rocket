../Small84/Queue_113.sv