../Small21/AXI4Buffer_2.sv