../Full11/head_40x6.sv