../Small12/CoherenceManagerWrapper.sv