../Medium41/TLXbar.sv