../Small81/Repeater_1.sv