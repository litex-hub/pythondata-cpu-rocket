../Small21/TLMonitor_22.sv