../Small11/Queue_2.sv