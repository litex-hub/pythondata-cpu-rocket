../Small21/Queue_35.sv