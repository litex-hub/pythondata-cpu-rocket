../Small22/CLINT.sv