../Medium81/ClockSinkDomain.sv