../Small12/Repeater_1.sv