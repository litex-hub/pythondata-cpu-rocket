../Small21/IntXbar_3.sv