../Small21/TLInterconnectCoupler_5.sv