../Medium28/SystemBus.sv