../Small82/CLINT.sv