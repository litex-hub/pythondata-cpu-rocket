../Small12/Queue_87.sv