../Small41/TLBuffer_5.sv