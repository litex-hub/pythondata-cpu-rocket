../Small24/AXI4Fragmenter_1.sv