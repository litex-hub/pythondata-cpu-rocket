../Small11/TLDebugModule.sv