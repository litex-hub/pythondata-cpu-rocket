../Small42/TLMonitor_50.sv