../Small41/TLAsyncCrossingSource.sv