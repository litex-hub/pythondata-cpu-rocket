../Full11/head_2x4.sv