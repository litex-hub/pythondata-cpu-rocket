../Small21/TLMonitor_31.sv