../Small41/TLMonitor_17.sv