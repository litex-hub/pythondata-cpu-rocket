../Small24/MemoryBus.sv