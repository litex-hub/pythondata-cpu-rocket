../Medium84/TilePRCIDomain.sv