../Small22/TLInterconnectCoupler_2.sv