../Small42/TLBroadcastTracker.sv