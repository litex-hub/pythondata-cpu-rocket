../Small42/TLMonitor_25.sv