../Small11/TLDebugModuleInner.sv