../Small81/BroadcastFilter.sv