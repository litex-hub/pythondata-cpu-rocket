../Small82/TLBroadcastTracker_1.sv