../Full11/CSRFile.sv