../Medium21/Queue_90.sv