../Small12/TLMonitor_14.sv