../Small11/Queue_21.sv