../Medium81/IntSyncCrossingSource_57.sv