../Medium41/TLMonitor_29.sv