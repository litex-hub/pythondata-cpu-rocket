../Small41/Queue_47.sv