../Small12/TLFIFOFixer_2.sv