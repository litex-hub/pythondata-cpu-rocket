../Small41/TLDebugModuleInnerAsync.sv