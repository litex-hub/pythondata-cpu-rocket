../Small82/Repeater_2.sv