../Small11/TLInterconnectCoupler_10.sv