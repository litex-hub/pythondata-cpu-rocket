../Small41/TLMonitor_22.sv