../Small11/ram_2x72.sv