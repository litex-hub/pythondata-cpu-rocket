../Small18/TLMonitor_23.sv