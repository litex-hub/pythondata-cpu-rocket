../Small11/AXI4IdIndexer.sv