../Small88/TLFIFOFixer_4.sv