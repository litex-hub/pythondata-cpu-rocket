../Small82/TLBroadcast.sv