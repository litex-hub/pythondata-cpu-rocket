../Small28/Queue_101.sv