../Small81/BundleBridgeNexus_78.sv