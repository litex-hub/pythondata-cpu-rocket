../Small41/Queue_101.sv