../Small22/TLToAXI4_1.sv