../Small21/TLMonitor_32.sv