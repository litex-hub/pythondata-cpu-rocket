../Medium81/ExampleRocketSystem.sv