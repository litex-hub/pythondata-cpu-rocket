../Medium12/ExampleRocketSystem.sv