../Full11/PMPChecker_2.sv