../Small48/TLBroadcastTracker_3.sv