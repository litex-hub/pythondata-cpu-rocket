../Small41/TLDebugModuleOuter.sv