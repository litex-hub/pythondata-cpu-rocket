../Small22/AXI4Buffer_2.sv