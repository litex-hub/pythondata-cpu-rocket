../Small81/AXI4UserYanker_2.sv