../Full11/OptimizationBarrier_37.sv