../Small11/Queue_36.sv