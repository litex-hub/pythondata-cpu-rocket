../Small44/Queue_101.sv