../Small41/TLXbar_16.sv