../Linux11/MulAddRecFNToRaw_postMul_1.sv