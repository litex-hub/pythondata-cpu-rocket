../Medium24/ExampleRocketSystem.sv