../Small12/TLMonitor_13.sv