../Small42/TLBuffer_4.sv