../Small41/Queue_54.sv