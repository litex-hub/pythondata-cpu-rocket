../Full11/SinkE.sv