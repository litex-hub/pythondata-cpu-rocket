../Linux41/RocketTile.sv