../Linux11/PTW.sv