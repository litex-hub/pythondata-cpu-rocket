../Medium84/ExampleRocketSystem.sv