../Full11/ICache.sv