../Small21/TLXbar_12.sv