../Small88/BankBinder.sv