../Small11/rf_31x64.sv