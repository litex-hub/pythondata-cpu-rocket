../Small18/TLToAXI4_1.sv