../Small82/TLMonitor_18.sv