../Small44/Queue_99.sv