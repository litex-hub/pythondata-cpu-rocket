../Small81/Queue_5.sv