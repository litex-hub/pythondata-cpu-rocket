../Small12/TLMonitor_33.sv