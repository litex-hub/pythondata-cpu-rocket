../Small14/ProbePicker.sv