../Small24/TLMonitor_21.sv