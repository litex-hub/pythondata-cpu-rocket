../Small12/TLMonitor_9.sv