../Small22/TLMonitor_32.sv