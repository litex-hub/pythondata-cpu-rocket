../Small21/Queue_44.sv