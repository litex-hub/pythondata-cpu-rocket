../Small11/ram_2x124.sv