../Small14/MemoryBus.sv