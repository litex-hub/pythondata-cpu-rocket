../Small41/TLMonitor_41.sv