../Small12/Queue_93.sv