../Small11/ram_2x71.sv