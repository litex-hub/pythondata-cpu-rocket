../Small24/AXI4UserYanker_2.sv