../Small42/TLMonitor_22.sv