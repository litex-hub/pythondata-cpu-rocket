../Small12/TLAtomicAutomata_1.sv