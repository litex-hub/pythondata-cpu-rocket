../Small41/Queue_64.sv