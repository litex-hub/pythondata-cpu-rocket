../Small12/TLDebugModuleInner.sv