../Small11/AXI4Buffer_2.sv