../Small81/TLMonitor_29.sv