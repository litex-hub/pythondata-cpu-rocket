../Small48/TLBroadcastTracker.sv