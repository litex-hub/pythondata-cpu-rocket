../Small44/Queue_107.sv