../Small41/TLFIFOFixer_2.sv