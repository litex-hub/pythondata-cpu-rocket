../Small11/SimAXIMem.sv