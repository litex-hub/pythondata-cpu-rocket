../Small11/AsyncQueueSink.sv