../Small42/TLDebugModuleOuter.sv