../Small22/TLToAXI4.sv