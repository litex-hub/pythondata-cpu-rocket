../Small42/AXI4Xbar.sv