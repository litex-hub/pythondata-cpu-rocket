../Small41/Queue_107.sv