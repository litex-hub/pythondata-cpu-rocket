../Small12/Repeater.sv