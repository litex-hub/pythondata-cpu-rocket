../Small81/AXI4Buffer_1.sv