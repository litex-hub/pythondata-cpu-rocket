../Small81/Rocket.sv