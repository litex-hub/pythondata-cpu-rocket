../Small21/TLBroadcastTracker_2.sv