../Full21/CoherenceManagerWrapper.sv