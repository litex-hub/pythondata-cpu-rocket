../Small44/TLInterconnectCoupler_18.sv