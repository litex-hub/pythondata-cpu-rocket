../Small18/Queue_74.sv