../Small81/Queue_164.sv