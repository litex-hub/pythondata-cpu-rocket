../Small42/Queue_142.sv