../Small81/TLMonitor_61.sv