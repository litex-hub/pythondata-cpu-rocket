../Linux81/Rocket.sv