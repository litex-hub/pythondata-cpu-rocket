../Small22/TLMonitor_36.sv