../Small11/Queue_38.sv