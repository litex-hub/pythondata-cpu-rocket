../Small22/TLMonitor_21.sv