../Small84/Repeater.sv