../Small22/TLMonitor_13.sv