../Small44/TLBroadcastTracker_2.sv