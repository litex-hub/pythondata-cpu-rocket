../Small41/TLInterconnectCoupler_7.sv