../Linux11/BTB.sv