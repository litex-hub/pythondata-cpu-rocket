../Small84/TLXbar.sv