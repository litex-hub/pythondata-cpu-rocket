../Small12/AXI4Fragmenter_1.sv