../Small21/AXI4ToTL.sv