../Small21/Queue_88.sv