../Small41/TLXbar_5.sv