../Small84/AXI4IdIndexer_2.sv