../Small81/ClockSinkDomain_1.sv