../Medium11/TLMonitor_25.sv