../Small41/TLMonitor_12.sv