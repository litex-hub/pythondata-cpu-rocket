../Small82/BankBinder.sv