../Small82/TLFragmenter_3.sv