../Small82/TLBroadcastTracker_3.sv