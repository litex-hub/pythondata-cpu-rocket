../Small11/TLInterconnectCoupler_8.sv