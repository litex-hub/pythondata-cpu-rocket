../Small11/TLMonitor_12.sv