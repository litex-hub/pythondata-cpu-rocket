../Small81/Queue_73.sv