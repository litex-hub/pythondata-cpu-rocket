../Small82/TLMonitor_26.sv