../Small12/TLMonitor_6.sv