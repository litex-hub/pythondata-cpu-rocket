../Small21/TLMonitor_23.sv