../Small18/TLMonitor_19.sv