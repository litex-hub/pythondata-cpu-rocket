../Small21/TLMonitor_20.sv