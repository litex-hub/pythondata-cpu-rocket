../Small22/TLMonitor_25.sv