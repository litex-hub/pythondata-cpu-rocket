../Small11/AXI4Buffer_1.sv