../Small28/TLMonitor_23.sv