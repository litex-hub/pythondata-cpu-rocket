../Medium11/TLPLIC.sv