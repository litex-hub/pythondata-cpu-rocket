../Medium21/TLMonitor_4.sv