../Linux11/data_arrays_512x128.sv