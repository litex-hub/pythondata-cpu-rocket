../Small11/Queue_23.sv