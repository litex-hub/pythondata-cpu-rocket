../Small12/TLDebugModuleOuter.sv