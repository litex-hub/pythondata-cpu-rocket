../Small22/TLMonitor_23.sv