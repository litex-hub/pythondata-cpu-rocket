../Small44/TLMonitor_29.sv