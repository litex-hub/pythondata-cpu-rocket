../Small21/Queue_97.sv