../Small42/TLMonitor_49.sv