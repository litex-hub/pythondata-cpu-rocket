../Small21/TLInterconnectCoupler_6.sv