../Small11/TLFIFOFixer_4.sv