../Small12/mem_134217728x128.sv