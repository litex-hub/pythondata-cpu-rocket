../Small42/TLXbar_8.sv