../Medium84/TLXbar.sv