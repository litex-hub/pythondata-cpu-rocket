../Full11/ram_12x109.sv