../Small41/TLMonitor_14.sv