../Small48/TLBroadcast.sv