../Small41/Queue_33.sv