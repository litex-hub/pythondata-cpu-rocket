../Small81/TLInterconnectCoupler_12.sv