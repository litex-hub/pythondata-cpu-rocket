../Small41/BankBinder.sv