../Medium41/RocketTile.sv