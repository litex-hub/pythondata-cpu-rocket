../Small12/TLMonitor_15.sv