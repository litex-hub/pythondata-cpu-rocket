../Medium21/TLXbar_8.sv