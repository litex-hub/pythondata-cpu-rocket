../Small82/AXI4Fragmenter_1.sv