../Full14/TilePRCIDomain.sv