../Small42/TLMonitor_11.sv