../Small41/TLMonitor_48.sv