../Small11/RVCExpander.sv