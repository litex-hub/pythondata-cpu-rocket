../Small11/data_arrays_512x32.sv