../Small22/TLMonitor_38.sv