../Small41/TLBroadcastTracker_3.sv