../Small11/Queue_91.sv