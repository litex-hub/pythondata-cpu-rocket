../Small48/TLBroadcastTracker_1.sv