../Full12/DCache.sv