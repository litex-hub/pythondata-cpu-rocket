../Small84/TLBroadcastTracker_1.sv