../Small28/AXI4UserYanker_2.sv