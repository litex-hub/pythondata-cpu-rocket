../Small12/ram_2x136.sv