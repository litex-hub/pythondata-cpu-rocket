../Linux11/FPU.sv