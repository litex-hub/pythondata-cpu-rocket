../Small82/AXI4Buffer_1.sv