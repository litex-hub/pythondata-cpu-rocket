../Small12/TLFragmenter_2.sv