../Small22/TLMonitor_11.sv