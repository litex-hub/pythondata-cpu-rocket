../Small81/Queue_61.sv