../Small22/TLMonitor_41.sv