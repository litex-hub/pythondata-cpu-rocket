../Small11/IntSyncAsyncCrossingSink.sv