../Linux41/CSRFile.sv