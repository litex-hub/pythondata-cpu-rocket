../Small41/TLMonitor_19.sv