../Medium41/Queue_105.sv