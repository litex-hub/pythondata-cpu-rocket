../Small82/TLMonitor_28.sv