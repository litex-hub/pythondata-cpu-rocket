../Small82/TLBroadcastTracker.sv