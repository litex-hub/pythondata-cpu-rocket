../Small11/TLMonitor_22.sv