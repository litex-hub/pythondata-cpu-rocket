../Small24/TLWidthWidget_2.sv