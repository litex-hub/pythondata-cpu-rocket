../Small11/PTW.sv