../Linux11/FPUDecoder.sv