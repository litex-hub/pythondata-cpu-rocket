../Small12/TLMonitor_5.sv