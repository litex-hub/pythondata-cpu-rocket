../Medium11/ram_2x109.sv