../Small11/Queue_35.sv