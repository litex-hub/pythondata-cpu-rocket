../Small11/IntSyncCrossingSource_4.sv