../Small44/TLMonitor_26.sv