../Small11/ClockSinkDomain.sv