../Small11/ram_2x73.sv