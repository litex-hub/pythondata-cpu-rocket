../Small81/RocketTile.sv