../Full11/TLMonitor.sv