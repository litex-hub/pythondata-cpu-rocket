../Small41/TLMonitor_21.sv