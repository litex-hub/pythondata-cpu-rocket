../Small21/TLInterconnectCoupler_9.sv