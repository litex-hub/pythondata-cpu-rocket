../Medium48/SystemBus.sv