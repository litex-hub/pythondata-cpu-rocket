../Small28/TLMonitor_24.sv