../Small11/TLDebugModuleOuter.sv