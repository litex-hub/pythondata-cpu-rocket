../Small28/TLMonitor_22.sv