../Small18/TLBroadcastTracker_1.sv