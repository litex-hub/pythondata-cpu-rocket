../Small81/AXI4Xbar_1.sv