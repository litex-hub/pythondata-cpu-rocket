../Small18/AXI4Xbar.sv