../Linux11/MulAddRecFNToRaw_preMul.sv