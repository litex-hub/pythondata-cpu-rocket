../Small11/ram_8x14.sv