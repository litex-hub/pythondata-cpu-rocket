../Small82/TLMonitor_35.sv