../Linux11/FPUFMAPipe.sv