../Small14/mem_67108864x256.sv