../Small12/Repeater_2.sv