../Linux11/RoundAnyRawFNToRecFN.sv