../Full11/data_33x45.sv