../Small81/TLMonitor_19.sv