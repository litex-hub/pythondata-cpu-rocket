../Small22/TLPLIC.sv