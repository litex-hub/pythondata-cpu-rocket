../Small41/IntXbar_5.sv