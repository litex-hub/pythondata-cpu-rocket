../Small14/TLMonitor_21.sv