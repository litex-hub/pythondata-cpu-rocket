../Small11/SimpleClockGroupSource.sv