../Small12/TLMonitor_24.sv