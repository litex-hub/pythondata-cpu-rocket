../Small41/TLFragmenter_1.sv