../Small44/TLXbar.sv