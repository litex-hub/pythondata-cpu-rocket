../Linux11/DivSqrtRecFNToRaw_small.sv