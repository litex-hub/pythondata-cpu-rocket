../Small21/Queue_91.sv