../Medium11/SystemBus.sv