../Small41/TLMonitor_50.sv