../Small22/Queue_81.sv