../Small12/TLBroadcastTracker.sv