../Full81/CSRFile.sv