../Small48/TLWidthWidget_2.sv