../Full11/ListBuffer.sv