../Small18/BankBinder.sv