../Small11/TLToAXI4_1.sv