../Small81/TLMonitor_63.sv