../Small11/Queue_22.sv