../Small81/TLAsyncCrossingSource.sv