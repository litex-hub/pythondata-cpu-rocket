../Small21/TLFragmenter_3.sv