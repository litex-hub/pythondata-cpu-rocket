../Small21/TLBroadcastTracker_1.sv