../Small11/TLMonitor_14.sv