../Medium22/TLPLIC.sv