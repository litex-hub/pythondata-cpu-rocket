../Small11/TLMonitor_18.sv