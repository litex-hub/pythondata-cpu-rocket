../Small41/TLFragmenter_3.sv