../Medium41/TLXbar_8.sv