../Linux11/table_512x1.sv