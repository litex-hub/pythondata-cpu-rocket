../Small11/TLMonitor_7.sv