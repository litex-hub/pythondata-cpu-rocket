../Full11/AXI4IdIndexer_2.sv