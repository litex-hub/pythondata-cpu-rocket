../Small11/ram_2x60.sv