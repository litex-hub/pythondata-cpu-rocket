../Full11/data_40x73.sv