../Small41/Queue_65.sv