../Small41/AsyncQueueSink_2.sv