../Small11/BreakpointUnit.sv