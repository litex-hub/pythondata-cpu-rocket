../Small88/CoherenceManagerWrapper.sv