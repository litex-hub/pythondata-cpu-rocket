../Small22/TLFragmenter_2.sv