../Medium24/SystemBus.sv