../Small41/Queue_50.sv