../Medium22/ExampleRocketSystem.sv