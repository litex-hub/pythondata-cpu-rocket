../Small22/Repeater_1.sv