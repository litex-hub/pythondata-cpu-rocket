../Small21/Queue_30.sv