../Small11/Queue_88.sv