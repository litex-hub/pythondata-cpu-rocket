../Small11/AXI4UserYanker.sv