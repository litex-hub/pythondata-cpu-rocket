../Small84/Repeater_1.sv