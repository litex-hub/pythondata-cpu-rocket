../Small82/TLError_1.sv