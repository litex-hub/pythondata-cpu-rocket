../Small42/TLMonitor_24.sv