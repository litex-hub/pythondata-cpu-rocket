../Small41/TLError_1.sv