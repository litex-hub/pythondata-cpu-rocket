../Small21/Queue_41.sv