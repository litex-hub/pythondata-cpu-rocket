../Medium81/TLMonitor_37.sv