../Medium18/SystemBus.sv