../Small42/TLMonitor_17.sv