../Small82/TLXbar_5.sv