../Small22/Queue_107.sv