../Small12/TLMonitor_7.sv