../Small12/TLFragmenter_1.sv