../Small21/Queue_43.sv