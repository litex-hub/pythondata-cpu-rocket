../Small41/TLMonitor_49.sv