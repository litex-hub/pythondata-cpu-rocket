../Small12/TLMonitor_19.sv