../Medium81/TLXbar.sv