../Small11/ram_2x79.sv