../Small81/AXI4Deinterleaver.sv