../Small21/TLMonitor_12.sv