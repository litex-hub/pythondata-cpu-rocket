../Small11/AXI4Buffer.sv