../Small11/TLBuffer_4.sv