../Full24/TilePRCIDomain.sv