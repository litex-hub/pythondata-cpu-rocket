../Small14/TLBroadcastTracker_1.sv