../Small21/AXI4Buffer_1.sv