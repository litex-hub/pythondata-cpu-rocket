../Medium81/Queue_111.sv