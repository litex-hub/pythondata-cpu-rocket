../Small12/TLMonitor_35.sv