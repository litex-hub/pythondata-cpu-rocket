../Small14/SimAXIMem.sv