../Small11/Queue_4.sv