../Small11/Queue_80.sv