../Small41/TLMonitor_20.sv