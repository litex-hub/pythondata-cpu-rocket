../Small48/TLFIFOFixer_4.sv