../Small82/TLBuffer_5.sv