../Small11/IntSyncSyncCrossingSink_1.sv