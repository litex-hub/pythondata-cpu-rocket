../Small18/Queue_87.sv