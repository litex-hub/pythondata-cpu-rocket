../Medium11/DCache.sv