../Small11/Queue_20.sv