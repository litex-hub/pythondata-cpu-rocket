../Linux81/FPU.sv