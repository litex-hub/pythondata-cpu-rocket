../Small41/ClockSinkDomain.sv