../Small11/DebugCustomXbar.sv