../Small11/IntSyncCrossingSource_1.sv