../Small12/TLMonitor_8.sv