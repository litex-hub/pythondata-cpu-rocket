../Small41/IntSyncCrossingSource_17.sv