../Small41/TLInterconnectCoupler_8.sv