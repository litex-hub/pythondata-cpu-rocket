../Medium82/TLFIFOFixer.sv