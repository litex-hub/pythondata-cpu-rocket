../Full11/next_33x6.sv