../Medium41/TLFIFOFixer.sv