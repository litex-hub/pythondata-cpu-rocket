../Small14/AXI4Fragmenter_1.sv