../Small41/TLDebugModule.sv