../Small84/MemoryBus.sv