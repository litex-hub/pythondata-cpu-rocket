../Small14/ram_2x288.sv