../Small48/Queue_99.sv