../Small11/Queue_90.sv