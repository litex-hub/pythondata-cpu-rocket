../Medium42/TLMonitor_30.sv