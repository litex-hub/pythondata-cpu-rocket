../Small41/AXI4Fragmenter.sv