../Small11/TLInterconnectCoupler_12.sv