../Small41/AXI4Fragmenter_2.sv