../Small42/TLError.sv