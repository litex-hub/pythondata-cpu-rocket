../Small42/TLMonitor_14.sv