../Full11/tail_40x6.sv