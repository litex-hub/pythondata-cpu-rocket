../Small11/TLBroadcastTracker_1.sv