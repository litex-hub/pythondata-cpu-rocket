../Linux11/tag_array_64x88.sv