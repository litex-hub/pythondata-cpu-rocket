../Small81/TLMonitor_25.sv