../Small12/Queue_72.sv