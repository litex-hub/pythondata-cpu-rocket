../Small42/TLMonitor_51.sv