../Small42/MemoryBus.sv