../Small81/Queue_107.sv