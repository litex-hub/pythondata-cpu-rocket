../Small21/IntSyncCrossingSource_9.sv