../Small21/TLMonitor_38.sv