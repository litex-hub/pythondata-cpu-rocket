../Medium28/ExampleRocketSystem.sv