../Small18/TLMonitor_22.sv