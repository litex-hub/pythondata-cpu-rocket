../Small41/Queue_55.sv