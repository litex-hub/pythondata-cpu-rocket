../Small41/AXI4ToTL.sv