../Small21/Queue_37.sv