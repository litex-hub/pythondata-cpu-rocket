../Small82/Repeater_5.sv