../Small11/TLMonitor_30.sv