../Small21/TLMonitor_39.sv