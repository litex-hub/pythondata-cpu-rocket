../Medium41/TLMonitor_31.sv