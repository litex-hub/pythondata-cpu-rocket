../Medium84/SystemBus.sv