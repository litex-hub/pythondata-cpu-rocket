../Linux11/Rocket.sv