../Small48/ProbePicker.sv