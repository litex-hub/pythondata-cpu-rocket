../Small44/Queue_132.sv