../Small84/Queue_161.sv