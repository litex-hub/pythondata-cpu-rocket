../Small42/TLMonitor_18.sv