../Medium41/CSRFile.sv