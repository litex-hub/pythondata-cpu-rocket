../Small11/TLError.sv