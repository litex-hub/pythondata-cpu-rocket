../Linux11/RocketTile.sv