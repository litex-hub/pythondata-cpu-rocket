../Small24/TLXbar.sv