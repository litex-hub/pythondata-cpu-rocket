../Small82/TLToAXI4_1.sv