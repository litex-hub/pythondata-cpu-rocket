../Small88/Queue_155.sv