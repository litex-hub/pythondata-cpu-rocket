../Full11/IBuf.sv