../Medium21/IntSyncCrossingSource_15.sv