../Small11/ResetSynchronizerShiftReg_w1_d3_i0.sv