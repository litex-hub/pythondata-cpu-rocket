../Small12/TLBroadcastTracker_1.sv