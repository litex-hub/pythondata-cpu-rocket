../Linux11/ICache.sv