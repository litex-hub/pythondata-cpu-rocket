../Small82/TLMonitor_33.sv