../Linux11/MulAddRecFNPipe_1.sv