../Small11/ProbePicker.sv