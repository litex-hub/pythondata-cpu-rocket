../Small11/TLMonitor_29.sv