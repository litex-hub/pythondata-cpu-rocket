../Small21/AXI4Fragmenter.sv