../Medium88/ExampleRocketSystem.sv