../Small21/TLError.sv