../Small24/TLMonitor_4.sv