../Small14/TLWidthWidget_2.sv