../Small48/Queue_101.sv