../Medium11/TLMonitor_23.sv