../Small11/Repeater_2.sv