../Small12/AXI4Buffer_1.sv