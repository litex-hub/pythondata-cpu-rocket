../Small11/TLMonitor_15.sv