../Small12/ram_2x145.sv