../Small22/AXI4Fragmenter_1.sv