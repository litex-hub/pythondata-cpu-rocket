../Small11/Queue_32.sv