../Small82/TLFragmenter_2.sv