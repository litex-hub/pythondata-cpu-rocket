../Small11/TLMonitor_2.sv