../Small14/TLBroadcastTracker_3.sv