../Medium18/ExampleRocketSystem.sv