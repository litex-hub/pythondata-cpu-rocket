../Small14/TLMonitor_3.sv