../Small42/TLXbar_5.sv