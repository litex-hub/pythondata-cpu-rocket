../Small84/Queue_107.sv