../Small11/Rocket.sv