../Small81/TLDebugModuleInner.sv