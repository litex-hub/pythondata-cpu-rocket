../Full11/tail_2x4.sv