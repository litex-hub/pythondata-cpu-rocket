../Small22/TLBroadcastTracker_1.sv