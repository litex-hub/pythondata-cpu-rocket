../Small11/TLMonitor_5.sv