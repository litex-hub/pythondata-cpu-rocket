../Small11/TLMonitor_13.sv