../Medium11/Arbiter.sv