../Small42/TLBusBypassBar.sv