../Medium41/ExampleRocketSystem.sv