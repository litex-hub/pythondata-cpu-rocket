../Small22/TLMonitor_6.sv