../Small11/FixedClockBroadcast_3.sv