../Small82/AXI4IdIndexer_2.sv