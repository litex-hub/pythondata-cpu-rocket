../Small24/TLBroadcastTracker.sv