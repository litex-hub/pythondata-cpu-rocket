../Small22/TLXbar_5.sv