../Small82/TLMonitor_32.sv