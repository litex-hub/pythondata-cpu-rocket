../Small28/TLFIFOFixer_4.sv