../Small18/MemoryBus.sv