../Small81/TLInterconnectCoupler_14.sv