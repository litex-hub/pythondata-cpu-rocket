../Small82/Queue_105.sv