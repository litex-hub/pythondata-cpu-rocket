../Full11/PMPChecker.sv