../Small41/MemoryBus.sv