../Small41/TLAtomicAutomata_1.sv