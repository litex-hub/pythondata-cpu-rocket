../Medium21/TLMonitor_26.sv