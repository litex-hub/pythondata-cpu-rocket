../Small81/TLFIFOFixer_2.sv