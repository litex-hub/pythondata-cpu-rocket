../Small41/Queue_132.sv