../Small14/TLFIFOFixer.sv