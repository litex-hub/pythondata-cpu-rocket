../Small82/TLError.sv