../Small41/Queue_125.sv