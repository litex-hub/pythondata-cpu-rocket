../Small11/CLINT.sv