../Small22/TLMonitor_24.sv