../Small12/TLMonitor_25.sv