../Small21/AXI4UserYanker_2.sv