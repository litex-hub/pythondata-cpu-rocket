../Small81/Queue_169.sv