../Full41/CSRFile.sv