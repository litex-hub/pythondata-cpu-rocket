../Full11/ram_sink_2x3.sv