../Small22/TLMonitor_15.sv