../Linux41/FPU.sv