../Medium21/TilePRCIDomain.sv