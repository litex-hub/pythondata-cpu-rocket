../Small41/TLMonitor_24.sv