../Small82/TLInterconnectCoupler_2.sv