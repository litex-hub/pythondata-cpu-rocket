../Small18/ram_2x520.sv