../Small81/TLBuffer_2.sv