../Small11/Queue_6.sv