../Small81/AXI4ToTL.sv