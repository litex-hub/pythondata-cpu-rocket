../Small11/ram_2x102.sv