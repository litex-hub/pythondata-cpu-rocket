../Small42/TLMonitor_23.sv