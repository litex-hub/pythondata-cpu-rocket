../Small11/ClockCrossingReg_w15.sv