../Small11/TLMonitor_27.sv