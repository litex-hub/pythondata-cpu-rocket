../Full11/PTW.sv