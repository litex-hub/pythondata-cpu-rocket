../Small44/TLMonitor_27.sv