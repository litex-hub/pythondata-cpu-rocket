../Small12/TLFragmenter.sv