../Full11/OptimizationBarrier_36.sv