../Small81/TLMonitor_18.sv