../Small21/Queue_7.sv