../Small12/TLMonitor_20.sv