../Small82/TLMonitor_65.sv