../Small82/TLToAXI4.sv