../Small21/TLMonitor_36.sv