../Small18/ram_2x577.sv