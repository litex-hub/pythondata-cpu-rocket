../Small11/ClockCrossingReg_w43.sv