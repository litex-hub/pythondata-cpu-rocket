../Small81/TLFragmenter.sv