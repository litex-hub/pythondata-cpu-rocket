../Small22/TLMonitor_18.sv