../Small82/TLMonitor_20.sv