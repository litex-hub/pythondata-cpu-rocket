../Small81/Queue_59.sv