../Small82/TLMonitor_25.sv