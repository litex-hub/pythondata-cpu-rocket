../Small42/TLMonitor_29.sv