../Medium81/TLMonitor_10.sv