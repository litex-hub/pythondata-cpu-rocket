../Small22/AXI4UserYanker_2.sv