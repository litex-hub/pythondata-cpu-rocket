../Small81/TLMonitor_32.sv