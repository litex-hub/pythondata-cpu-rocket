../Small18/ProbePicker.sv