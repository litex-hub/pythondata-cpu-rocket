../Small11/Queue_74.sv