../Small18/TLInterconnectCoupler_12.sv