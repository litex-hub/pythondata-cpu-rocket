../Small24/Queue_104.sv