../Small14/AXI4Xbar.sv