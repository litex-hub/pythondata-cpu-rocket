../Small21/TLXbar_5.sv