../Small82/MemoryBus.sv