../Small11/TLBuffer_5.sv