../Linux11/FPUFMAPipe_1.sv