../Small12/BankBinder.sv