../Small88/Queue_158.sv