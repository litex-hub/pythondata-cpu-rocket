../Small41/FixedClockBroadcast.sv