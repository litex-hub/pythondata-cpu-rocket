../Medium88/SystemBus.sv