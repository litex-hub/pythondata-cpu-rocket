../Small22/TLMonitor_19.sv