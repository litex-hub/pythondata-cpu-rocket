../Small81/TLInterconnectCoupler_15.sv