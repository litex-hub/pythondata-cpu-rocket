../Small41/AXI4Xbar_1.sv