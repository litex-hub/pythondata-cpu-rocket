../Small41/BundleBridgeNexus_42.sv