../Small18/Queue_72.sv