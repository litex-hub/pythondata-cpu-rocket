../Small44/TLFIFOFixer_4.sv