../Medium81/TLMonitor_39.sv