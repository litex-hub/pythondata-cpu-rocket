../Medium81/RocketTile.sv