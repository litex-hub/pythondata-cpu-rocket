../Full81/Rocket.sv