../Small81/FixedClockBroadcast.sv