../Medium21/TLMonitor_1.sv