../Small81/IntSyncCrossingSource_49.sv