../Small21/TLBusBypassBar.sv