../Small84/TLMonitor_33.sv