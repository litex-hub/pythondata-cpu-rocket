../Full11/Repeater_1.sv