../Medium42/TLMonitor_6.sv