../Small22/TLMonitor_8.sv