../Small11/ClockCrossingReg_w55.sv