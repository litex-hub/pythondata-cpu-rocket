../Small12/TLBusBypassBar.sv