../Medium11/ICache.sv