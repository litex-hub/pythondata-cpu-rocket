../Small21/Queue_100.sv