../Small81/TLDebugModuleOuter.sv