../Small42/TLError_1.sv