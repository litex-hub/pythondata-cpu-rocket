../Medium24/TLXbar.sv