../Small12/TLFragmenter_3.sv