../Small88/AXI4UserYanker_2.sv