../Small41/TLMonitor_23.sv