../Small18/TLInterconnectCoupler_2.sv