../Small28/CoherenceManagerWrapper.sv