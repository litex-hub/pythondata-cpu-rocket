../Small82/TLBusBypassBar.sv