../Small11/AXI4UserYanker_1.sv