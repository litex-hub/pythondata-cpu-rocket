../Small44/AXI4Buffer_1.sv