../Small48/TLBroadcastTracker_2.sv