../Medium11/ExampleRocketSystem.sv