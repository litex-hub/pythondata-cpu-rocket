../Small82/TLMonitor_24.sv