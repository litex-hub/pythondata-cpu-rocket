../Small41/TLMonitor_5.sv