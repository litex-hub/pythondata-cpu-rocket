../Small42/TLMonitor_10.sv