../Linux11/RoundAnyRawFNToRecFN_4.sv