../Small21/TLMonitor_3.sv