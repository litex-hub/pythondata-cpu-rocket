../Medium22/TLXbar_8.sv