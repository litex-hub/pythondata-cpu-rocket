../Medium42/TLFIFOFixer.sv