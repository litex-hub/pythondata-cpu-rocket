../Medium81/Rocket.sv