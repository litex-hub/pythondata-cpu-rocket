../Small11/Queue_84.sv