../Small22/MemoryBus.sv