../Small42/TLFIFOFixer_4.sv