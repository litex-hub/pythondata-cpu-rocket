../Small41/TLMonitor_10.sv