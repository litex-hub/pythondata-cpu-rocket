../Small84/TLMonitor_18.sv