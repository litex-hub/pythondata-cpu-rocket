../Small21/TLMonitor_19.sv