../Small11/MaxPeriodFibonacciLFSR.sv