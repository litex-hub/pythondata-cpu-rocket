../Small84/BankBinder.sv