../Small41/TLMonitor_15.sv