../Full11/Atomics.sv