../Small11/Queue_37.sv