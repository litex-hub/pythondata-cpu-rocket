../Small42/TLBroadcastTracker_1.sv