../Linux81/RocketTile.sv