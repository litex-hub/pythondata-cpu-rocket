../Full12/ICache.sv