../Small81/TLError.sv