../Small11/DCache.sv