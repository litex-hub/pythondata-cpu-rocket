../Small41/TLBroadcast.sv