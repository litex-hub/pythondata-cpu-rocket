../Linux11/data_arrays_0_512x256.sv