../Small82/TLInterconnectCoupler_26.sv