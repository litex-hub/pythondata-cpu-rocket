../Small81/IntSyncCrossingSource_33.sv