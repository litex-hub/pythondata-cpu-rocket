../Small11/Queue_86.sv