../Small22/Queue_101.sv