../Small41/TLBuffer_2.sv