../Small82/TLFIFOFixer_3.sv