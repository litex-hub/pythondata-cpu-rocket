../Small18/Queue_90.sv