../Small18/TLBroadcastTracker_3.sv