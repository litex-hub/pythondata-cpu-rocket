../Small41/TLInterconnectCoupler_18.sv