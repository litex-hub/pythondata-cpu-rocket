../Small11/Frontend.sv