../Medium11/TLMonitor_3.sv