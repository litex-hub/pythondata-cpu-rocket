../Small81/TLMonitor_20.sv