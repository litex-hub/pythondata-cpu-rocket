../Medium82/TLMonitor_40.sv