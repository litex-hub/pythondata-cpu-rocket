../Small11/TLToAXI4.sv