../Small14/TLBroadcastTracker_2.sv