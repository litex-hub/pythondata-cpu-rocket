../Small22/TLInterconnectCoupler_14.sv