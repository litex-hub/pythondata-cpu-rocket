../Small41/IntSyncCrossingSource_25.sv