../Medium21/TLMonitor_25.sv