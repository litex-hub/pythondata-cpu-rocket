../Medium21/TLBuffer_10.sv