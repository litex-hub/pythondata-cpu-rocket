../Medium12/TLFIFOFixer.sv