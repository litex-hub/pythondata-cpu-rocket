../Small41/TLMonitor_44.sv