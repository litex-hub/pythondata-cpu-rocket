../Small24/Queue_81.sv