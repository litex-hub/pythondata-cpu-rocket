../Small84/CoherenceManagerWrapper.sv