../Small41/TLBuffer_4.sv