../Small11/IntSyncCrossingSource_7.sv