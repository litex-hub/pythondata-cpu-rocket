../Small11/Queue_1.sv