../Small84/TLFIFOFixer_4.sv