../Medium81/SystemBus.sv