../Small41/Queue_53.sv