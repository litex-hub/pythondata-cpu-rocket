../Small81/ErrorDeviceWrapper.sv