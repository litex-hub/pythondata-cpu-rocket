../Small21/TLDebugModuleOuter.sv