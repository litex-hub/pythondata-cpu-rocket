../Small11/HellaCacheArbiter.sv