../Small21/Queue_36.sv