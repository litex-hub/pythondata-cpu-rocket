../Small21/Queue_29.sv