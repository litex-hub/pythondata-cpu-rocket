../Small11/AXI4Fragmenter_1.sv