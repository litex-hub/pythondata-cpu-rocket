../Small14/AXI4UserYanker_2.sv