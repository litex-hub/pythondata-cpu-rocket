../Small44/AXI4UserYanker_2.sv