../Small28/Queue_81.sv