../Small42/TLMonitor_21.sv