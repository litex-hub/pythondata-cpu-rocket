../Small11/AXI4RAM_1.sv