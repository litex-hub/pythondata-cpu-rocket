../Small44/TLBroadcastTracker_1.sv