../Small11/TLMonitor_4.sv