../Medium41/ClockSinkDomain.sv