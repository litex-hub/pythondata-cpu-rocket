../Small81/TLMonitor_26.sv