../Small81/Queue_55.sv