../Small42/TLAsyncCrossingSource.sv