../Small11/ram_8x72.sv