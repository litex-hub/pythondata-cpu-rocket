../Small41/TLError.sv