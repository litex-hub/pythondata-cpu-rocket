../Small41/TLBuffer_3.sv