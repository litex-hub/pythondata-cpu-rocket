../Small82/TLMonitor_36.sv