../Full11/tail_21x6.sv