../Medium11/TLB_1.sv