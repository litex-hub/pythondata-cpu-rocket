../Small82/TLFIFOFixer_4.sv