../Small11/MemoryBus.sv