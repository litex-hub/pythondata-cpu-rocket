../Small28/TLMonitor_21.sv