../Small21/Queue_32.sv