../Medium41/TilePRCIDomain.sv