../Full11/ListBuffer_1.sv