../Small11/TLROM.sv