../Small11/CoherenceManagerWrapper.sv