../Small88/Queue_161.sv