../Small21/TLFragmenter_1.sv