../Full11/Repeater_3.sv