../Full11/BTB.sv