../Small18/mem_33554432x512.sv