../Medium82/TLMonitor_10.sv