../Small11/Queue.sv