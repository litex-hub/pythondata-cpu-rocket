../Small18/AXI4IdIndexer_2.sv