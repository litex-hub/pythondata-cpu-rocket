../Small81/ram_16x16.sv