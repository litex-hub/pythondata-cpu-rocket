../Small84/TLMonitor_37.sv