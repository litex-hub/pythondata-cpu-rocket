../Small11/AXI4UserYanker_2.sv