../Medium81/TLFIFOFixer.sv