../Small18/TLBroadcast.sv