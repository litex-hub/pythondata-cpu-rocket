../Medium12/TLXbar.sv