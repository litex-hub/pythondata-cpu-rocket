../Small81/TLBroadcast.sv