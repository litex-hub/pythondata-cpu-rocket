../Small11/ICache.sv