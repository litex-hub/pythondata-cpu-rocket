../Medium11/TLXbar_8.sv