../Small81/Queue_112.sv