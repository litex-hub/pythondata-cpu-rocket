../Small82/TLDebugModuleInner.sv