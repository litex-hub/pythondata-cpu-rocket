../Small22/TLBroadcastTracker_2.sv