../Small21/Queue_115.sv