../Small48/BankBinder.sv