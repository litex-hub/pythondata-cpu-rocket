../Small21/TLBroadcastTracker_3.sv