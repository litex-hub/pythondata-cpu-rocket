../Small22/TLDebugModuleOuter.sv