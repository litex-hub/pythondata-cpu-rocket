../Small82/TLMonitor_66.sv