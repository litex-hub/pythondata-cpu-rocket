../Linux11/MulAddRecFNToRaw_postMul.sv