../Small42/TLFragmenter_2.sv