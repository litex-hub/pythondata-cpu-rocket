../Small88/TLMonitor_33.sv