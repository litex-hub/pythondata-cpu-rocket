../Small22/TLDebugModuleInner.sv