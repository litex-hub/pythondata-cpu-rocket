../Small41/Queue_59.sv