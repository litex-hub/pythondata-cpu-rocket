../Small21/Queue_47.sv