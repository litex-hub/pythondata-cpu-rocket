../Small81/Repeater.sv