../Small11/Queue_26.sv