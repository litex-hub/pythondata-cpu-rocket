../Small42/TLFragmenter.sv