../Small84/AXI4Xbar.sv