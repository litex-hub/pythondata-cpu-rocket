../Small81/Queue_53.sv