../Small41/Queue_143.sv