../Small21/TLAtomicAutomata_1.sv