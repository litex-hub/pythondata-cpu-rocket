../Small11/AMOALU.sv