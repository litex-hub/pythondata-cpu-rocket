../Small48/AXI4Fragmenter_1.sv