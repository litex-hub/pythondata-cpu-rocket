../Small42/Queue_129.sv