../Small42/AXI4Buffer_2.sv