../Small11/BroadcastFilter.sv