../Small84/TLWidthWidget_2.sv