../Medium42/TLXbar.sv