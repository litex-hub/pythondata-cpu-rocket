../Medium21/ExampleRocketSystem.sv