../Small11/AsyncResetSynchronizerPrimitiveShiftReg_d3_i0.sv