../Small21/TLAsyncCrossingSource.sv