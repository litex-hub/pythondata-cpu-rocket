../Small11/AsyncValidSync.sv