../Small81/TLMonitor_27.sv