../Small22/TLBroadcastTracker_3.sv