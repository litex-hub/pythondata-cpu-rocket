../Small24/Repeater_1.sv