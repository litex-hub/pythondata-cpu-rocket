../Small21/TLInterconnectCoupler_14.sv