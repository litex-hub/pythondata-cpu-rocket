../Small22/TLBuffer_5.sv