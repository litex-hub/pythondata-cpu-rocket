../Small48/TLMonitor_28.sv