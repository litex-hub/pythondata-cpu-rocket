../Small44/TLWidthWidget_2.sv