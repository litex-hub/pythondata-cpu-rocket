../Small28/TLMonitor_25.sv