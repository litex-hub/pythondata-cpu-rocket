../Small21/TLToAXI4_1.sv