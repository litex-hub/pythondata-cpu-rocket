../Medium11/BreakpointUnit.sv