../Small22/TLFIFOFixer_4.sv