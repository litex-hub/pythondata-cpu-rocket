../Medium44/ExampleRocketSystem.sv