../Small11/AXI4Deinterleaver.sv