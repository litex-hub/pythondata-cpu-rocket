../Small11/ShiftQueue.sv