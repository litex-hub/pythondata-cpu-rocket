../Small81/TLMonitor_69.sv