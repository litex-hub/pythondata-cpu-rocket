../Small81/TLBusBypassBar.sv