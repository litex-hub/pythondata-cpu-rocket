../Small14/TLMonitor_20.sv