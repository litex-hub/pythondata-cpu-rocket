../Medium21/SystemBus.sv