../Small11/ALU.sv