../Small81/TLBuffer_3.sv