../Small11/ErrorDeviceWrapper.sv