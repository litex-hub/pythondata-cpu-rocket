../Small42/TLROM.sv