../Small82/TLDebugModuleOuter.sv