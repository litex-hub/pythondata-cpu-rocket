../Small22/TLMonitor_34.sv