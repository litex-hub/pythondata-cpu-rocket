../Small81/Queue_152.sv