../Small41/Queue_61.sv