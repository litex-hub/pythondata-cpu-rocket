../Small11/TLMonitor_31.sv