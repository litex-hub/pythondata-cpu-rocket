../Medium42/TLPLIC.sv