../Medium41/IntSyncCrossingSource_29.sv