../Small11/ram_8x9.sv