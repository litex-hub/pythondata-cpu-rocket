../Small82/TLMonitor_31.sv