../Small12/TLMonitor_17.sv