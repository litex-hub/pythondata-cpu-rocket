../Medium82/TLMonitor_39.sv