../Small88/TLInterconnectCoupler_2.sv