../Small82/TLMonitor_22.sv