../Small12/TLMonitor_30.sv