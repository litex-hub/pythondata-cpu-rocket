../Small82/CoherenceManagerWrapper.sv