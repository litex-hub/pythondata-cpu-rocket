../Small12/TLError_1.sv