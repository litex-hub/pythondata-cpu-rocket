../Medium12/TLXbar_8.sv