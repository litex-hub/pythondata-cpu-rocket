../Small24/TLBuffer_10.sv