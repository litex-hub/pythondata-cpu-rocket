../Small22/TLBroadcast.sv