../Small11/AsyncQueueSource_1.sv