../Small42/TLBroadcast.sv