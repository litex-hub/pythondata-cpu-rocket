../Small14/ram_2x289.sv