../Small88/TLMonitor_35.sv