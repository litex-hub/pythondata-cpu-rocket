../Small41/Queue_126.sv