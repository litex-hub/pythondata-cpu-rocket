../Small82/TLMonitor_30.sv