../Full11/ram_2x80.sv