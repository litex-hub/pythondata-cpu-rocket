../Small41/TLFragmenter.sv