../Small42/TLWidthWidget_2.sv