../Small41/CLINT.sv