../Small44/AXI4Xbar.sv