../Small11/ram_2x62.sv