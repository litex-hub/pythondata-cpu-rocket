../Small21/TLBroadcast.sv