../Small28/Queue_104.sv