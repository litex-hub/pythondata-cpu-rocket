../Small42/TLMonitor_43.sv