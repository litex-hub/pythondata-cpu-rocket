../Small88/AXI4Buffer_1.sv