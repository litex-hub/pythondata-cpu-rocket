../Full42/RocketTile.sv