../Small21/ProbePicker.sv