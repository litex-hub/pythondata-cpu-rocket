../Medium22/TilePRCIDomain.sv