../Small82/TLMonitor_23.sv