../Small11/MulDiv.sv