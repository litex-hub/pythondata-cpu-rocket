../Small81/Queue_54.sv