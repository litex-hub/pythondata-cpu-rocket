../Small24/TLMonitor_24.sv