../Small48/TLMonitor_27.sv