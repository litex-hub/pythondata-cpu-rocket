../Small82/TLBuffer_2.sv