../Small22/TLFIFOFixer_3.sv