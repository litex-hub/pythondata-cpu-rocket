../Small12/SimAXIMem.sv