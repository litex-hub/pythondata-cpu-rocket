../Small82/TLMonitor_21.sv