../Small18/TLWidthWidget_2.sv