../Small11/TLMonitor_20.sv