../Small81/AXI4Fragmenter.sv