../Small11/TLMonitor_17.sv