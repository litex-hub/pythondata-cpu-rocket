../Small81/Queue_56.sv