../Medium41/TLMonitor_30.sv