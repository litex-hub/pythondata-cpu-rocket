../Small24/TLFIFOFixer_4.sv