../Small12/TLMonitor_16.sv