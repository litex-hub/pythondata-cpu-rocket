../Small81/TLMonitor_66.sv