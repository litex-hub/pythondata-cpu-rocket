../Small14/TLInterconnectCoupler_12.sv