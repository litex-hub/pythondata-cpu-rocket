../Small12/Repeater_5.sv