../Small24/TLMonitor_25.sv