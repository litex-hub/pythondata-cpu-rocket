../Small44/TLMonitor_28.sv