../Small11/TLAsyncCrossingSink.sv