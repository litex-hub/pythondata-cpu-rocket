../Full21/TLMonitor_1.sv