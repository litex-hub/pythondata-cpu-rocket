../Small21/TLBuffer_2.sv