../Small81/Queue_115.sv