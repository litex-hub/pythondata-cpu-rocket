../Small81/TLMonitor_34.sv