../Small81/ram_8x82.sv