../Small41/AXI4UserYanker.sv