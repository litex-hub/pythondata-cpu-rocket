../Small21/TLBuffer_3.sv