../Small12/TLXbar_5.sv