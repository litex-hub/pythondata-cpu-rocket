../Small41/TLDebugModuleOuterAsync.sv