../Small21/AXI4Deinterleaver.sv