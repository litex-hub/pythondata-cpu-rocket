../Small12/TLMonitor_31.sv