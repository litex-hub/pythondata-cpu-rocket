../Small41/TLMonitor_47.sv