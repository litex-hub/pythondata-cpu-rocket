../Small11/SynchronizerShiftReg_w1_d3.sv