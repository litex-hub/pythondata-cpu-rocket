../Small81/TLBroadcastTracker_3.sv