../Medium42/TLBuffer_10.sv