../Small44/TLMonitor_6.sv