../Small11/Queue_101.sv