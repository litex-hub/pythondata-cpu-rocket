../Small48/AXI4Buffer_1.sv