../Small81/TLBroadcastTracker_1.sv