../Small82/TLMonitor_68.sv