../Small81/AsyncQueueSource_1.sv