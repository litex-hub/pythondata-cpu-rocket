../Small41/AXI4Deinterleaver.sv