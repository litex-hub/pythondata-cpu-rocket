../Small11/TLMonitor_19.sv