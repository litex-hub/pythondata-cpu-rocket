../Small41/TLDebugModuleInner.sv