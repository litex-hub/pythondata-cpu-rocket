../Medium22/TLMonitor_4.sv