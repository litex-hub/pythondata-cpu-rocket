../Small18/AXI4Fragmenter_1.sv