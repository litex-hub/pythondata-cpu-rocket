../Medium44/TLFIFOFixer.sv