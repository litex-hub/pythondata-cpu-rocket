../Small84/Queue_155.sv