../Small28/Repeater_1.sv