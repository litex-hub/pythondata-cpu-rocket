../Small11/ram_2x116.sv