../Small21/AXI4UserYanker_1.sv