../Medium41/SystemBus.sv